** Generated for: hspiceD
** Generated on: Sep 14 17:59:54 2014
** Design library name: dummy_4_bit
** Design cell name: test_OAI21
** Design view name: schematic
.GLOBAL vdd! _gnet0 vss!
.PARAM cap=0.663f vdd=1 v_low=0 buff_vdd=vdd v_hig=vdd


.TRAN 100e-12 1e-6 START=0.0

.OP

.TEMP 25
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
+    post=1
.PROBE TRAN V(a) V(b1) V(b2) V(a_in) V(b1_in) V(b2_in) V(output) V(Vpower)
.INCLUDE "/ad/eng/users/b/o/bobzhou/Desktop/571/hw3/tech_files/45nm_HP.pm"

** Library name: NangateOpenCellLibrary
** Cell name: OAI21_X2
** View name: schematic
.subckt OAI21_X2 a b1 b2 zn
m_i_2_0 vss! a net_0 vss! NMOS_VTL L=50e-9 W=415e-9
m_i_2_1 net_0 a vss! vss! NMOS_VTL L=50e-9 W=415e-9
m_i_1__m0 zn b2 net_0 vss! NMOS_VTL L=50e-9 W=415e-9
m_i_1__m1 net_0 b2 zn vss! NMOS_VTL L=50e-9 W=415e-9
m_i_0__m0 net_0 b1 zn vss! NMOS_VTL L=50e-9 W=415e-9
m_i_0__m1 zn b1 net_0 vss! NMOS_VTL L=50e-9 W=415e-9
m_i_3__m0 zn b1 net_1__m0_0 _gnet0 PMOS_VTL L=50e-9 W=630e-9
m_i_4__m0 net_1__m0_0 b2 _gnet0 _gnet0 PMOS_VTL L=50e-9 W=630e-9
m_i_3__m1 net_1__m1 b1 zn _gnet0 PMOS_VTL L=50e-9 W=630e-9
m_i_4__m1 _gnet0 b2 net_1__m1 _gnet0 PMOS_VTL L=50e-9 W=630e-9
m_i_5_0 zn a _gnet0 _gnet0 PMOS_VTL L=50e-9 W=630e-9
m_i_5_1 _gnet0 a zn _gnet0 PMOS_VTL L=50e-9 W=630e-9
.ends OAI21_X2
** End of subcircuit definition.

** Library name: equalized_logic
** Cell name: buffer4test
** View name: schematic
.subckt buffer4test buff_vdd buff_vss input output inh_bulk_n inh_bulk_p
m1 output net14 buff_vdd inh_bulk_p pmos_vtl L=50e-9 W=1.26e-6
m3 net14 input buff_vdd inh_bulk_p pmos_vtl L=50e-9 W=1.26e-6
m0 output net14 buff_vss inh_bulk_n nmos_vtl L=50e-9 W=830e-9
m9 net14 input buff_vss inh_bulk_n nmos_vtl L=50e-9 W=830e-9
.ends buffer4test
** End of subcircuit definition.

** Library name: dummy_4_bit
** Cell name: test_OAI21
** View name: schematic
xi15 a_in b1_in b2_in output OAI21_X2
f0 vpower 0 CCCS v3  1 M=1
v10 buff_vss 0 DC=0
v8 buff_vdd 0 DC=buff_vdd
v6 vss! 0 DC=0
v3 _gnet0 0 DC=vdd
xi18 buff_vdd buff_vss b2 b2_in 0 vdd! buffer4test
xi17 buff_vdd buff_vss b1 b1_in 0 vdd! buffer4test
xi16 buff_vdd buff_vss a a_in 0 vdd! buffer4test
c10 vpower 0 1e-12 IC=0
c0 output 0 663e-18
v4 b2 0 PWL
+ 1.000000000e-12 V_hig
+ 1.000000000e-09 V_hig
+ 1.001000000e-09 V_hig
+ 1.100000000e-09 V_hig
+ 1.101000000e-09 V_hig
+ 1.200000000e-09 V_hig
+ 1.201000000e-09 V_hig
+ 1.300000000e-09 V_hig
+ 1.301000000e-09 V_hig
+ 1.400000000e-09 V_hig
+ 1.401000000e-09 V_hig
+ 1.500000000e-09 V_hig
+ 1.501000000e-09 V_hig
+ 1.600000000e-09 V_hig
+ 1.601000000e-09 V_hig
+ 1.700000000e-09 V_hig
+ 1.701000000e-09 V_hig
+ 1.800000000e-09 V_hig
+ 1.801000000e-09 V_hig
+ 1.900000000e-09 V_hig
+ 1.901000000e-09 V_hig
+ 2.000000000e-09 V_hig
+ 2.001000000e-09 V_hig
+ 2.100000000e-09 V_hig
+ 2.101000000e-09 V_hig
+ 2.200000000e-09 V_hig
+ 2.201000000e-09 V_hig
+ 2.300000000e-09 V_hig
+ 2.301000000e-09 V_hig
+ 2.400000000e-09 V_hig
+ 2.401000000e-09 V_hig
+ 2.500000000e-09 V_hig
+ 2.501000000e-09 V_hig
+ 2.600000000e-09 V_hig
+ 2.601000000e-09 V_hig
+ 2.700000000e-09 V_hig
+ 2.701000000e-09 V_hig
+ 2.800000000e-09 V_hig
+ 2.801000000e-09 V_hig
+ 2.900000000e-09 V_hig
+ 2.901000000e-09 V_low
+ 3.000000000e-09 V_low
+ 3.001000000e-09 V_low
+ 3.100000000e-09 V_low
+ 3.101000000e-09 V_low
+ 3.200000000e-09 V_low
+ 3.201000000e-09 V_low
+ 3.300000000e-09 V_low
+ 3.301000000e-09 V_low
+ 3.400000000e-09 V_low
+ 3.401000000e-09 V_low
+ 3.500000000e-09 V_low
+ 3.501000000e-09 V_low
+ 3.600000000e-09 V_low
+ 3.601000000e-09 V_low
+ 3.700000000e-09 V_low
+ 3.701000000e-09 V_low
+ 3.800000000e-09 V_low
+ 3.801000000e-09 V_low
+ 3.900000000e-09 V_low
+ 3.901000000e-09 V_low
+ 4.000000000e-09 V_low
+ 4.001000000e-09 V_low
+ 4.100000000e-09 V_low
+ 4.101000000e-09 V_low
+ 4.200000000e-09 V_low
+ 4.201000000e-09 V_low
+ 4.300000000e-09 V_low
+ 4.301000000e-09 V_low
+ 4.400000000e-09 V_low
+ 4.401000000e-09 V_low
+ 4.500000000e-09 V_low
+ 4.501000000e-09 V_low
+ 4.600000000e-09 V_low
+ 4.601000000e-09 V_low
+ 4.700000000e-09 V_low
+ 4.701000000e-09 V_low
+ 4.800000000e-09 V_low
+ 4.801000000e-09 V_low
+ 4.900000000e-09 V_low
+ 4.901000000e-09 V_hig
+ 5.000000000e-09 V_hig
+ 5.001000000e-09 V_hig
+ 5.100000000e-09 V_hig
+ 5.101000000e-09 V_hig
+ 5.200000000e-09 V_hig
+ 5.201000000e-09 V_hig
+ 5.300000000e-09 V_hig
+ 5.301000000e-09 V_hig
+ 5.400000000e-09 V_hig
+ 5.401000000e-09 V_hig
+ 5.500000000e-09 V_hig
+ 5.501000000e-09 V_hig
+ 5.600000000e-09 V_hig
+ 5.601000000e-09 V_hig
+ 5.700000000e-09 V_hig
+ 5.701000000e-09 V_hig
+ 5.800000000e-09 V_hig
+ 5.801000000e-09 V_hig
+ 5.900000000e-09 V_hig
+ 5.901000000e-09 V_low
+ 6.000000000e-09 V_low
+ 6.001000000e-09 V_low
+ 6.100000000e-09 V_low
+ 6.101000000e-09 V_low
+ 6.200000000e-09 V_low
+ 6.201000000e-09 V_low
+ 6.300000000e-09 V_low
+ 6.301000000e-09 V_low
+ 6.400000000e-09 V_low
+ 6.401000000e-09 V_low
+ 6.500000000e-09 V_low
+ 6.501000000e-09 V_low
+ 6.600000000e-09 V_low
+ 6.601000000e-09 V_low
+ 6.700000000e-09 V_low
+ 6.701000000e-09 V_low
+ 6.800000000e-09 V_low
+ 6.801000000e-09 V_low
+ 6.900000000e-09 V_low
+ 6.901000000e-09 V_hig
+ 7.000000000e-09 V_hig
+ 7.001000000e-09 V_hig
+ 7.100000000e-09 V_hig
+ 7.101000000e-09 V_hig
+ 7.200000000e-09 V_hig
+ 7.201000000e-09 V_hig
+ 7.300000000e-09 V_hig
+ 7.301000000e-09 V_hig
+ 7.400000000e-09 V_hig
+ 7.401000000e-09 V_hig
+ 7.500000000e-09 V_hig
+ 7.501000000e-09 V_hig
+ 7.600000000e-09 V_hig
+ 7.601000000e-09 V_hig
+ 7.700000000e-09 V_hig
+ 7.701000000e-09 V_hig
+ 7.800000000e-09 V_hig
+ 7.801000000e-09 V_hig
+ 7.900000000e-09 V_hig
+ 7.901000000e-09 V_low
+ 8.000000000e-09 V_low
+ 8.001000000e-09 V_low
+ 8.100000000e-09 V_low
+ 8.101000000e-09 V_low
+ 8.200000000e-09 V_low
+ 8.201000000e-09 V_low
+ 8.300000000e-09 V_low
+ 8.301000000e-09 V_low
+ 8.400000000e-09 V_low
+ 8.401000000e-09 V_low
+ 8.500000000e-09 V_low
+ 8.501000000e-09 V_low
+ 8.600000000e-09 V_low
+ 8.601000000e-09 V_low
+ 8.700000000e-09 V_low
+ 8.701000000e-09 V_low
+ 8.800000000e-09 V_low
+ 8.801000000e-09 V_low
+ 8.900000000e-09 V_low
+ 8.901000000e-09 V_low
+ 9.000000000e-09 V_low
+ 9.001000000e-09 V_low
+ 9.100000000e-09 V_low
+ 9.101000000e-09 V_low
+ 9.200000000e-09 V_low
+ 9.201000000e-09 V_low
+ 9.300000000e-09 V_low
+ 9.301000000e-09 V_low
+ 9.400000000e-09 V_low
+ 9.401000000e-09 V_low
+ 9.500000000e-09 V_low
+ 9.501000000e-09 V_low
+ 9.600000000e-09 V_low
+ 9.601000000e-09 V_low
+ 9.700000000e-09 V_low
+ 9.701000000e-09 V_low
+ 9.800000000e-09 V_low
+ 9.801000000e-09 V_low
+ 9.900000000e-09 V_low
+ 9.901000000e-09 V_hig
+ 1.000000000e-08 V_hig
+ 1.000100000e-08 V_hig
+ 1.010000000e-08 V_hig
+ 1.010100000e-08 V_hig
+ 1.020000000e-08 V_hig
+ 1.020100000e-08 V_hig
+ 1.030000000e-08 V_hig
+ 1.030100000e-08 V_hig
+ 1.040000000e-08 V_hig
+ 1.040100000e-08 V_hig
+ 1.050000000e-08 V_hig
+ 1.050100000e-08 V_hig
+ 1.060000000e-08 V_hig
+ 1.060100000e-08 V_hig
+ 1.070000000e-08 V_hig
+ 1.070100000e-08 V_hig
+ 1.080000000e-08 V_hig
+ 1.080100000e-08 V_hig
+ 1.090000000e-08 V_hig
+ 1.090100000e-08 V_low
+ 1.100000000e-08 V_low
+ 1.100100000e-08 V_low
+ 1.110000000e-08 V_low
+ 1.110100000e-08 V_low
+ 1.120000000e-08 V_low
+ 1.120100000e-08 V_low
+ 1.130000000e-08 V_low
+ 1.130100000e-08 V_low
+ 1.140000000e-08 V_low
+ 1.140100000e-08 V_low
+ 1.150000000e-08 V_low
+ 1.150100000e-08 V_low
+ 1.160000000e-08 V_low
+ 1.160100000e-08 V_low
+ 1.170000000e-08 V_low
+ 1.170100000e-08 V_low
+ 1.180000000e-08 V_low
+ 1.180100000e-08 V_low
+ 1.190000000e-08 V_low
+ 1.190100000e-08 V_hig
+ 1.200000000e-08 V_hig
+ 1.200100000e-08 V_hig
+ 1.210000000e-08 V_hig
+ 1.210100000e-08 V_hig
+ 1.220000000e-08 V_hig
+ 1.220100000e-08 V_hig
+ 1.230000000e-08 V_hig
+ 1.230100000e-08 V_hig
+ 1.240000000e-08 V_hig
+ 1.240100000e-08 V_hig
+ 1.250000000e-08 V_hig
+ 1.250100000e-08 V_hig
+ 1.260000000e-08 V_hig
+ 1.260100000e-08 V_hig
+ 1.270000000e-08 V_hig
+ 1.270100000e-08 V_hig
+ 1.280000000e-08 V_hig
+ 1.280100000e-08 V_hig
+ 1.290000000e-08 V_hig
+ 1.290100000e-08 V_low
+ 1.300000000e-08 V_low
+ 1.300100000e-08 V_low
+ 1.310000000e-08 V_low
+ 1.310100000e-08 V_low
+ 1.320000000e-08 V_low
+ 1.320100000e-08 V_low
+ 1.330000000e-08 V_low
+ 1.330100000e-08 V_low
+ 1.340000000e-08 V_low
+ 1.340100000e-08 V_low
+ 1.350000000e-08 V_low
+ 1.350100000e-08 V_low
+ 1.360000000e-08 V_low
+ 1.360100000e-08 V_low
+ 1.370000000e-08 V_low
+ 1.370100000e-08 V_low
+ 1.380000000e-08 V_low
+ 1.380100000e-08 V_low
+ 1.390000000e-08 V_low
+ 1.390100000e-08 V_hig
+ 1.400000000e-08 V_hig
+ 1.400100000e-08 V_hig
+ 1.410000000e-08 V_hig
+ 1.410100000e-08 V_hig
+ 1.420000000e-08 V_hig
+ 1.420100000e-08 V_hig
+ 1.430000000e-08 V_hig
+ 1.430100000e-08 V_hig
+ 1.440000000e-08 V_hig
+ 1.440100000e-08 V_hig
+ 1.450000000e-08 V_hig
+ 1.450100000e-08 V_hig
+ 1.460000000e-08 V_hig
+ 1.460100000e-08 V_hig
+ 1.470000000e-08 V_hig
+ 1.470100000e-08 V_hig
+ 1.480000000e-08 V_hig
+ 1.480100000e-08 V_hig
+ 1.490000000e-08 V_hig
+ 1.490100000e-08 V_hig
+ 1.500000000e-08 V_hig
+ 1.500100000e-08 V_hig
+ 1.510000000e-08 V_hig
+ 1.510100000e-08 V_hig
+ 1.520000000e-08 V_hig
+ 1.520100000e-08 V_hig
+ 1.530000000e-08 V_hig
+ 1.530100000e-08 V_hig
+ 1.540000000e-08 V_hig
+ 1.540100000e-08 V_hig
+ 1.550000000e-08 V_hig
+ 1.550100000e-08 V_hig
+ 1.560000000e-08 V_hig
+ 1.560100000e-08 V_hig
+ 1.570000000e-08 V_hig
+ 1.570100000e-08 V_hig
+ 1.580000000e-08 V_hig
+ 1.580100000e-08 V_hig
+ 1.590000000e-08 V_hig
+ 1.590100000e-08 V_hig
+ 1.600000000e-08 V_hig
+ 1.600100000e-08 V_hig
+ 1.610000000e-08 V_hig
+ 1.610100000e-08 V_hig
+ 1.620000000e-08 V_hig
+ 1.620100000e-08 V_hig
+ 1.630000000e-08 V_hig
+ 1.630100000e-08 V_hig
+ 1.640000000e-08 V_hig
+ 1.640100000e-08 V_hig
+ 1.650000000e-08 V_hig
+ 1.650100000e-08 V_hig
+ 1.660000000e-08 V_hig
+ 1.660100000e-08 V_hig
+ 1.670000000e-08 V_hig
+ 1.670100000e-08 V_hig
+ 1.680000000e-08 V_hig
+ 1.680100000e-08 V_hig
+ 1.690000000e-08 V_hig
+ 1.690100000e-08 V_hig
+ 1.700000000e-08 V_hig
+ 1.700100000e-08 V_hig
+ 1.710000000e-08 V_hig
+ 1.710100000e-08 V_hig
+ 1.720000000e-08 V_hig
+ 1.720100000e-08 V_hig
+ 1.730000000e-08 V_hig
+ 1.730100000e-08 V_hig
+ 1.740000000e-08 V_hig
+ 1.740100000e-08 V_hig
+ 1.750000000e-08 V_hig
+ 1.750100000e-08 V_hig
+ 1.760000000e-08 V_hig
+ 1.760100000e-08 V_hig
+ 1.770000000e-08 V_hig
+ 1.770100000e-08 V_hig
+ 1.780000000e-08 V_hig
+ 1.780100000e-08 V_hig
+ 1.790000000e-08 V_hig
+ 1.790100000e-08 V_hig
+ 1.800000000e-08 V_hig
+ 1.800100000e-08 V_hig
+ 1.810000000e-08 V_hig
+ 1.810100000e-08 V_hig
+ 1.820000000e-08 V_hig
+ 1.820100000e-08 V_hig
+ 1.830000000e-08 V_hig
+ 1.830100000e-08 V_hig
+ 1.840000000e-08 V_hig
+ 1.840100000e-08 V_hig
+ 1.850000000e-08 V_hig
+ 1.850100000e-08 V_hig
+ 1.860000000e-08 V_hig
+ 1.860100000e-08 V_hig
+ 1.870000000e-08 V_hig
+ 1.870100000e-08 V_hig
+ 1.880000000e-08 V_hig
+ 1.880100000e-08 V_hig
+ 1.890000000e-08 V_hig
+ 1.890100000e-08 V_low
+ 1.900000000e-08 V_low
+ 1.900100000e-08 V_low
+ 1.910000000e-08 V_low
+ 1.910100000e-08 V_low
+ 1.920000000e-08 V_low
+ 1.920100000e-08 V_low
+ 1.930000000e-08 V_low
+ 1.930100000e-08 V_low
+ 1.940000000e-08 V_low
+ 1.940100000e-08 V_low
+ 1.950000000e-08 V_low
+ 1.950100000e-08 V_low
+ 1.960000000e-08 V_low
+ 1.960100000e-08 V_low
+ 1.970000000e-08 V_low
+ 1.970100000e-08 V_low
+ 1.980000000e-08 V_low
+ 1.980100000e-08 V_low
+ 1.990000000e-08 V_low
+ 1.990100000e-08 V_hig
+ 2.000000000e-08 V_hig
+ 2.000100000e-08 V_hig
+ 2.010000000e-08 V_hig
+ 2.010100000e-08 V_hig
+ 2.020000000e-08 V_hig
+ 2.020100000e-08 V_hig
+ 2.030000000e-08 V_hig
+ 2.030100000e-08 V_hig
+ 2.040000000e-08 V_hig
+ 2.040100000e-08 V_hig
+ 2.050000000e-08 V_hig
+ 2.050100000e-08 V_hig
+ 2.060000000e-08 V_hig
+ 2.060100000e-08 V_hig
+ 2.070000000e-08 V_hig
+ 2.070100000e-08 V_hig
+ 2.080000000e-08 V_hig
+ 2.080100000e-08 V_hig
+ 2.090000000e-08 V_hig
+ 2.090100000e-08 V_hig
+ 2.100000000e-08 V_hig
+ 2.100100000e-08 V_hig
+ 2.110000000e-08 V_hig
+ 2.110100000e-08 V_hig
+ 2.120000000e-08 V_hig
+ 2.120100000e-08 V_hig
+ 2.130000000e-08 V_hig
+ 2.130100000e-08 V_hig
+ 2.140000000e-08 V_hig
+ 2.140100000e-08 V_hig
+ 2.150000000e-08 V_hig
+ 2.150100000e-08 V_hig
+ 2.160000000e-08 V_hig
+ 2.160100000e-08 V_hig
+ 2.170000000e-08 V_hig
+ 2.170100000e-08 V_hig
+ 2.180000000e-08 V_hig
+ 2.180100000e-08 V_hig
+ 2.190000000e-08 V_hig
+ 2.190100000e-08 V_low
+ 2.200000000e-08 V_low
+ 2.200100000e-08 V_low
+ 2.210000000e-08 V_low
+ 2.210100000e-08 V_low
+ 2.220000000e-08 V_low
+ 2.220100000e-08 V_low
+ 2.230000000e-08 V_low
+ 2.230100000e-08 V_low
+ 2.240000000e-08 V_low
+ 2.240100000e-08 V_low
+ 2.250000000e-08 V_low
+ 2.250100000e-08 V_low
+ 2.260000000e-08 V_low
+ 2.260100000e-08 V_low
+ 2.270000000e-08 V_low
+ 2.270100000e-08 V_low
+ 2.280000000e-08 V_low
+ 2.280100000e-08 V_low
+ 2.290000000e-08 V_low
+ 2.290100000e-08 V_hig
+ 2.300000000e-08 V_hig
+ 2.300100000e-08 V_hig
+ 2.310000000e-08 V_hig
+ 2.310100000e-08 V_hig
+ 2.320000000e-08 V_hig
+ 2.320100000e-08 V_hig
+ 2.330000000e-08 V_hig
+ 2.330100000e-08 V_hig
+ 2.340000000e-08 V_hig
+ 2.340100000e-08 V_hig
+ 2.350000000e-08 V_hig
+ 2.350100000e-08 V_hig
+ 2.360000000e-08 V_hig
+ 2.360100000e-08 V_hig
+ 2.370000000e-08 V_hig
+ 2.370100000e-08 V_hig
+ 2.380000000e-08 V_hig
+ 2.380100000e-08 V_hig
+ 2.390000000e-08 V_hig
+ 2.390100000e-08 V_hig
+ 2.400000000e-08 V_hig
+ 2.400100000e-08 V_hig
+ 2.410000000e-08 V_hig
+ 2.410100000e-08 V_hig
+ 2.420000000e-08 V_hig
+ 2.420100000e-08 V_hig
+ 2.430000000e-08 V_hig
+ 2.430100000e-08 V_hig
+ 2.440000000e-08 V_hig
+ 2.440100000e-08 V_hig
+ 2.450000000e-08 V_hig
+ 2.450100000e-08 V_hig
+ 2.460000000e-08 V_hig
+ 2.460100000e-08 V_hig
+ 2.470000000e-08 V_hig
+ 2.470100000e-08 V_hig
+ 2.480000000e-08 V_hig
+ 2.480100000e-08 V_hig
+ 2.490000000e-08 V_hig
+ 2.490100000e-08 V_low
+ 2.500000000e-08 V_low
+ 2.500100000e-08 V_low
+ 2.510000000e-08 V_low
+ 2.510100000e-08 V_low
+ 2.520000000e-08 V_low
+ 2.520100000e-08 V_low
+ 2.530000000e-08 V_low
+ 2.530100000e-08 V_low
+ 2.540000000e-08 V_low
+ 2.540100000e-08 V_low
+ 2.550000000e-08 V_low
+ 2.550100000e-08 V_low
+ 2.560000000e-08 V_low
+ 2.560100000e-08 V_low
+ 2.570000000e-08 V_low
+ 2.570100000e-08 V_low
+ 2.580000000e-08 V_low
+ 2.580100000e-08 V_low
+ 2.590000000e-08 V_low
+ 2.590100000e-08 V_low
+ 2.600000000e-08 V_low
+ 2.600100000e-08 V_low
+ 2.610000000e-08 V_low
+ 2.610100000e-08 V_low
+ 2.620000000e-08 V_low
+ 2.620100000e-08 V_low
+ 2.630000000e-08 V_low
+ 2.630100000e-08 V_low
+ 2.640000000e-08 V_low
+ 2.640100000e-08 V_low
+ 2.650000000e-08 V_low
+ 2.650100000e-08 V_low
+ 2.660000000e-08 V_low
+ 2.660100000e-08 V_low
+ 2.670000000e-08 V_low
+ 2.670100000e-08 V_low
+ 2.680000000e-08 V_low
+ 2.680100000e-08 V_low
+ 2.690000000e-08 V_low
+ 2.690100000e-08 V_hig
+ 2.700000000e-08 V_hig
+ 2.700100000e-08 V_hig
+ 2.710000000e-08 V_hig
+ 2.710100000e-08 V_hig
+ 2.720000000e-08 V_hig
+ 2.720100000e-08 V_hig
+ 2.730000000e-08 V_hig
+ 2.730100000e-08 V_hig
+ 2.740000000e-08 V_hig
+ 2.740100000e-08 V_hig
+ 2.750000000e-08 V_hig
+ 2.750100000e-08 V_hig
+ 2.760000000e-08 V_hig
+ 2.760100000e-08 V_hig
+ 2.770000000e-08 V_hig
+ 2.770100000e-08 V_hig
+ 2.780000000e-08 V_hig
+ 2.780100000e-08 V_hig
+ 2.790000000e-08 V_hig
+ 2.790100000e-08 V_low
+ 2.800000000e-08 V_low
+ 2.800100000e-08 V_low
+ 2.810000000e-08 V_low
+ 2.810100000e-08 V_low
+ 2.820000000e-08 V_low
+ 2.820100000e-08 V_low
+ 2.830000000e-08 V_low
+ 2.830100000e-08 V_low
+ 2.840000000e-08 V_low
+ 2.840100000e-08 V_low
+ 2.850000000e-08 V_low
+ 2.850100000e-08 V_low
+ 2.860000000e-08 V_low
+ 2.860100000e-08 V_low
+ 2.870000000e-08 V_low
+ 2.870100000e-08 V_low
+ 2.880000000e-08 V_low
+ 2.880100000e-08 V_low
+ 2.890000000e-08 V_low
+ 2.890100000e-08 V_low
+ 2.900000000e-08 V_low
+ 2.900100000e-08 V_low
+ 2.910000000e-08 V_low
+ 2.910100000e-08 V_low
+ 2.920000000e-08 V_low
+ 2.920100000e-08 V_low
+ 2.930000000e-08 V_low
+ 2.930100000e-08 V_low
+ 2.940000000e-08 V_low
+ 2.940100000e-08 V_low
+ 2.950000000e-08 V_low
+ 2.950100000e-08 V_low
+ 2.960000000e-08 V_low
+ 2.960100000e-08 V_low
+ 2.970000000e-08 V_low
+ 2.970100000e-08 V_low
+ 2.980000000e-08 V_low
+ 2.980100000e-08 V_low
+ 2.990000000e-08 V_low
+ 2.990100000e-08 V_low
+ 3.000000000e-08 V_low
+ 3.000100000e-08 V_low
+ 3.010000000e-08 V_low
+ 3.010100000e-08 V_low
+ 3.020000000e-08 V_low
+ 3.020100000e-08 V_low
+ 3.030000000e-08 V_low
+ 3.030100000e-08 V_low
+ 3.040000000e-08 V_low
+ 3.040100000e-08 V_low
+ 3.050000000e-08 V_low
+ 3.050100000e-08 V_low
+ 3.060000000e-08 V_low
+ 3.060100000e-08 V_low
+ 3.070000000e-08 V_low
+ 3.070100000e-08 V_low
+ 3.080000000e-08 V_low
+ 3.080100000e-08 V_low
+ 3.090000000e-08 V_low
+ 3.090100000e-08 V_hig
+ 3.100000000e-08 V_hig
+ 3.100100000e-08 V_hig
+ 3.110000000e-08 V_hig
+ 3.110100000e-08 V_hig
+ 3.120000000e-08 V_hig
+ 3.120100000e-08 V_hig
+ 3.130000000e-08 V_hig
+ 3.130100000e-08 V_hig
+ 3.140000000e-08 V_hig
+ 3.140100000e-08 V_hig
+ 3.150000000e-08 V_hig
+ 3.150100000e-08 V_hig
+ 3.160000000e-08 V_hig
+ 3.160100000e-08 V_hig
+ 3.170000000e-08 V_hig
+ 3.170100000e-08 V_hig
+ 3.180000000e-08 V_hig
+ 3.180100000e-08 V_hig
+ 3.190000000e-08 V_hig
+ 3.190100000e-08 V_hig
+ 3.200000000e-08 V_hig
+ 3.200100000e-08 V_hig
+ 3.210000000e-08 V_hig
+ 3.210100000e-08 V_hig
+ 3.220000000e-08 V_hig
+ 3.220100000e-08 V_hig
+ 3.230000000e-08 V_hig
+ 3.230100000e-08 V_hig
+ 3.240000000e-08 V_hig
+ 3.240100000e-08 V_hig
+ 3.250000000e-08 V_hig
+ 3.250100000e-08 V_hig
+ 3.260000000e-08 V_hig
+ 3.260100000e-08 V_hig
+ 3.270000000e-08 V_hig
+ 3.270100000e-08 V_hig
+ 3.280000000e-08 V_hig
+ 3.280100000e-08 V_hig
+ 3.290000000e-08 V_hig
+ 3.290100000e-08 V_low
+ 3.300000000e-08 V_low
+ 3.300100000e-08 V_low
+ 3.310000000e-08 V_low
+ 3.310100000e-08 V_low
+ 3.320000000e-08 V_low
+ 3.320100000e-08 V_low
+ 3.330000000e-08 V_low
+ 3.330100000e-08 V_low
+ 3.340000000e-08 V_low
+ 3.340100000e-08 V_low
+ 3.350000000e-08 V_low
+ 3.350100000e-08 V_low
+ 3.360000000e-08 V_low
+ 3.360100000e-08 V_low
+ 3.370000000e-08 V_low
+ 3.370100000e-08 V_low
+ 3.380000000e-08 V_low
+ 3.380100000e-08 V_low
+ 3.390000000e-08 V_low
+ 3.390100000e-08 V_low
+ 3.400000000e-08 V_low
+ 3.400100000e-08 V_low
+ 3.410000000e-08 V_low
+ 3.410100000e-08 V_low
+ 3.420000000e-08 V_low
+ 3.420100000e-08 V_low
+ 3.430000000e-08 V_low
+ 3.430100000e-08 V_low
+ 3.440000000e-08 V_low
+ 3.440100000e-08 V_low
+ 3.450000000e-08 V_low
+ 3.450100000e-08 V_low
+ 3.460000000e-08 V_low
+ 3.460100000e-08 V_low
+ 3.470000000e-08 V_low
+ 3.470100000e-08 V_low
+ 3.480000000e-08 V_low
+ 3.480100000e-08 V_low
+ 3.490000000e-08 V_low
+ 3.490100000e-08 V_hig
+ 3.500000000e-08 V_hig
+ 3.500100000e-08 V_hig
+ 3.510000000e-08 V_hig
+ 3.510100000e-08 V_hig
+ 3.520000000e-08 V_hig
+ 3.520100000e-08 V_hig
+ 3.530000000e-08 V_hig
+ 3.530100000e-08 V_hig
+ 3.540000000e-08 V_hig
+ 3.540100000e-08 V_hig
+ 3.550000000e-08 V_hig
+ 3.550100000e-08 V_hig
+ 3.560000000e-08 V_hig
+ 3.560100000e-08 V_hig
+ 3.570000000e-08 V_hig
+ 3.570100000e-08 V_hig
+ 3.580000000e-08 V_hig
+ 3.580100000e-08 V_hig
+ 3.590000000e-08 V_hig
+ 3.590100000e-08 V_low
+ 3.600000000e-08 V_low
+ 3.600100000e-08 V_low
+ 3.610000000e-08 V_low
+ 3.610100000e-08 V_low
+ 3.620000000e-08 V_low
+ 3.620100000e-08 V_low
+ 3.630000000e-08 V_low
+ 3.630100000e-08 V_low
+ 3.640000000e-08 V_low
+ 3.640100000e-08 V_low
+ 3.650000000e-08 V_low
+ 3.650100000e-08 V_low
+ 3.660000000e-08 V_low
+ 3.660100000e-08 V_low
+ 3.670000000e-08 V_low
+ 3.670100000e-08 V_low
+ 3.680000000e-08 V_low
+ 3.680100000e-08 V_low
+ 3.690000000e-08 V_low
+ 3.690100000e-08 V_low
+ 3.700000000e-08 V_low
+ 3.700100000e-08 V_low
+ 3.710000000e-08 V_low
+ 3.710100000e-08 V_low
+ 3.720000000e-08 V_low
+ 3.720100000e-08 V_low
+ 3.730000000e-08 V_low
+ 3.730100000e-08 V_low
+ 3.740000000e-08 V_low
+ 3.740100000e-08 V_low
+ 3.750000000e-08 V_low
+ 3.750100000e-08 V_low
+ 3.760000000e-08 V_low
+ 3.760100000e-08 V_low
+ 3.770000000e-08 V_low
+ 3.770100000e-08 V_low
+ 3.780000000e-08 V_low
+ 3.780100000e-08 V_low
+ 3.790000000e-08 V_low
+ 3.790100000e-08 V_hig
+ 3.800000000e-08 V_hig
+ 3.800100000e-08 V_hig
+ 3.810000000e-08 V_hig
+ 3.810100000e-08 V_hig
+ 3.820000000e-08 V_hig
+ 3.820100000e-08 V_hig
+ 3.830000000e-08 V_hig
+ 3.830100000e-08 V_hig
+ 3.840000000e-08 V_hig
+ 3.840100000e-08 V_hig
+ 3.850000000e-08 V_hig
+ 3.850100000e-08 V_hig
+ 3.860000000e-08 V_hig
+ 3.860100000e-08 V_hig
+ 3.870000000e-08 V_hig
+ 3.870100000e-08 V_hig
+ 3.880000000e-08 V_hig
+ 3.880100000e-08 V_hig
+ 3.890000000e-08 V_hig
+ 3.890100000e-08 V_low
+ 3.900000000e-08 V_low
+ 3.900100000e-08 V_low
+ 3.910000000e-08 V_low
+ 3.910100000e-08 V_low
+ 3.920000000e-08 V_low
+ 3.920100000e-08 V_low
+ 3.930000000e-08 V_low
+ 3.930100000e-08 V_low
+ 3.940000000e-08 V_low
+ 3.940100000e-08 V_low
+ 3.950000000e-08 V_low
+ 3.950100000e-08 V_low
+ 3.960000000e-08 V_low
+ 3.960100000e-08 V_low
+ 3.970000000e-08 V_low
+ 3.970100000e-08 V_low
+ 3.980000000e-08 V_low
+ 3.980100000e-08 V_low
+ 3.990000000e-08 V_low
+ 3.990100000e-08 V_hig
+ 4.000000000e-08 V_hig
+ 4.000100000e-08 V_hig
+ 4.010000000e-08 V_hig
+ 4.010100000e-08 V_hig
+ 4.020000000e-08 V_hig
+ 4.020100000e-08 V_hig
+ 4.030000000e-08 V_hig
+ 4.030100000e-08 V_hig
+ 4.040000000e-08 V_hig
+ 4.040100000e-08 V_hig
+ 4.050000000e-08 V_hig
+ 4.050100000e-08 V_hig
+ 4.060000000e-08 V_hig
+ 4.060100000e-08 V_hig
+ 4.070000000e-08 V_hig
+ 4.070100000e-08 V_hig
+ 4.080000000e-08 V_hig
+ 4.080100000e-08 V_hig
+ 4.090000000e-08 V_hig
+ 4.090100000e-08 V_hig
+ 4.100000000e-08 V_hig
+ 4.100100000e-08 V_hig
+ 4.110000000e-08 V_hig
+ 4.110100000e-08 V_hig
+ 4.120000000e-08 V_hig
+ 4.120100000e-08 V_hig
+ 4.130000000e-08 V_hig
+ 4.130100000e-08 V_hig
+ 4.140000000e-08 V_hig
+ 4.140100000e-08 V_hig
+ 4.150000000e-08 V_hig
+ 4.150100000e-08 V_hig
+ 4.160000000e-08 V_hig
+ 4.160100000e-08 V_hig
+ 4.170000000e-08 V_hig
+ 4.170100000e-08 V_hig
+ 4.180000000e-08 V_hig
+ 4.180100000e-08 V_hig
+ 4.190000000e-08 V_hig
+ 4.190100000e-08 V_low
+ 4.200000000e-08 V_low
+ 4.200100000e-08 V_low
+ 4.210000000e-08 V_low
+ 4.210100000e-08 V_low
+ 4.220000000e-08 V_low
+ 4.220100000e-08 V_low
+ 4.230000000e-08 V_low
+ 4.230100000e-08 V_low
+ 4.240000000e-08 V_low
+ 4.240100000e-08 V_low
+ 4.250000000e-08 V_low
+ 4.250100000e-08 V_low
+ 4.260000000e-08 V_low
+ 4.260100000e-08 V_low
+ 4.270000000e-08 V_low
+ 4.270100000e-08 V_low
+ 4.280000000e-08 V_low
+ 4.280100000e-08 V_low
+ 4.290000000e-08 V_low
+ 4.290100000e-08 V_hig
+ 4.300000000e-08 V_hig
+ 4.300100000e-08 V_hig
+ 4.310000000e-08 V_hig
+ 4.310100000e-08 V_hig
+ 4.320000000e-08 V_hig
+ 4.320100000e-08 V_hig
+ 4.330000000e-08 V_hig
+ 4.330100000e-08 V_hig
+ 4.340000000e-08 V_hig
+ 4.340100000e-08 V_hig
+ 4.350000000e-08 V_hig
+ 4.350100000e-08 V_hig
+ 4.360000000e-08 V_hig
+ 4.360100000e-08 V_hig
+ 4.370000000e-08 V_hig
+ 4.370100000e-08 V_hig
+ 4.380000000e-08 V_hig
+ 4.380100000e-08 V_hig
+ 4.390000000e-08 V_hig
+ 4.390100000e-08 V_hig
+ 4.400000000e-08 V_hig
+ 4.400100000e-08 V_hig
+ 4.410000000e-08 V_hig
+ 4.410100000e-08 V_hig
+ 4.420000000e-08 V_hig
+ 4.420100000e-08 V_hig
+ 4.430000000e-08 V_hig
+ 4.430100000e-08 V_hig
+ 4.440000000e-08 V_hig
+ 4.440100000e-08 V_hig
+ 4.450000000e-08 V_hig
+ 4.450100000e-08 V_hig
+ 4.460000000e-08 V_hig
+ 4.460100000e-08 V_hig
+ 4.470000000e-08 V_hig
+ 4.470100000e-08 V_hig
+ 4.480000000e-08 V_hig
+ 4.480100000e-08 V_hig
+ 4.490000000e-08 V_hig
+ 4.490100000e-08 V_hig
+ 4.500000000e-08 V_hig
+ 4.500100000e-08 V_hig
+ 4.510000000e-08 V_hig
+ 4.510100000e-08 V_hig
+ 4.520000000e-08 V_hig
+ 4.520100000e-08 V_hig
+ 4.530000000e-08 V_hig
+ 4.530100000e-08 V_hig
+ 4.540000000e-08 V_hig
+ 4.540100000e-08 V_hig
+ 4.550000000e-08 V_hig
+ 4.550100000e-08 V_hig
+ 4.560000000e-08 V_hig
+ 4.560100000e-08 V_hig
+ 4.570000000e-08 V_hig
+ 4.570100000e-08 V_hig
+ 4.580000000e-08 V_hig
+ 4.580100000e-08 V_hig
+ 4.590000000e-08 V_hig
+ 4.590100000e-08 V_low
+ 4.600000000e-08 V_low
+ 4.600100000e-08 V_low
+ 4.610000000e-08 V_low
+ 4.610100000e-08 V_low
+ 4.620000000e-08 V_low
+ 4.620100000e-08 V_low
+ 4.630000000e-08 V_low
+ 4.630100000e-08 V_low
+ 4.640000000e-08 V_low
+ 4.640100000e-08 V_low
+ 4.650000000e-08 V_low
+ 4.650100000e-08 V_low
+ 4.660000000e-08 V_low
+ 4.660100000e-08 V_low
+ 4.670000000e-08 V_low
+ 4.670100000e-08 V_low
+ 4.680000000e-08 V_low
+ 4.680100000e-08 V_low
+ 4.690000000e-08 V_low
+ 4.690100000e-08 V_hig
+ 4.700000000e-08 V_hig
+ 4.700100000e-08 V_hig
+ 4.710000000e-08 V_hig
+ 4.710100000e-08 V_hig
+ 4.720000000e-08 V_hig
+ 4.720100000e-08 V_hig
+ 4.730000000e-08 V_hig
+ 4.730100000e-08 V_hig
+ 4.740000000e-08 V_hig
+ 4.740100000e-08 V_hig
+ 4.750000000e-08 V_hig
+ 4.750100000e-08 V_hig
+ 4.760000000e-08 V_hig
+ 4.760100000e-08 V_hig
+ 4.770000000e-08 V_hig
+ 4.770100000e-08 V_hig
+ 4.780000000e-08 V_hig
+ 4.780100000e-08 V_hig
+ 4.790000000e-08 V_hig
+ 4.790100000e-08 V_low
+ 4.800000000e-08 V_low
+ 4.800100000e-08 V_low
+ 4.810000000e-08 V_low
+ 4.810100000e-08 V_low
+ 4.820000000e-08 V_low
+ 4.820100000e-08 V_low
+ 4.830000000e-08 V_low
+ 4.830100000e-08 V_low
+ 4.840000000e-08 V_low
+ 4.840100000e-08 V_low
+ 4.850000000e-08 V_low
+ 4.850100000e-08 V_low
+ 4.860000000e-08 V_low
+ 4.860100000e-08 V_low
+ 4.870000000e-08 V_low
+ 4.870100000e-08 V_low
+ 4.880000000e-08 V_low
+ 4.880100000e-08 V_low
+ 4.890000000e-08 V_low
+ 4.890100000e-08 V_low
+ 4.900000000e-08 V_low
+ 4.900100000e-08 V_low
+ 4.910000000e-08 V_low
+ 4.910100000e-08 V_low
+ 4.920000000e-08 V_low
+ 4.920100000e-08 V_low
+ 4.930000000e-08 V_low
+ 4.930100000e-08 V_low
+ 4.940000000e-08 V_low
+ 4.940100000e-08 V_low
+ 4.950000000e-08 V_low
+ 4.950100000e-08 V_low
+ 4.960000000e-08 V_low
+ 4.960100000e-08 V_low
+ 4.970000000e-08 V_low
+ 4.970100000e-08 V_low
+ 4.980000000e-08 V_low
+ 4.980100000e-08 V_low
+ 4.990000000e-08 V_low
+ 4.990100000e-08 V_hig
+ 5.000000000e-08 V_hig
+ 5.000100000e-08 V_hig
+ 5.010000000e-08 V_hig
+ 5.010100000e-08 V_hig
+ 5.020000000e-08 V_hig
+ 5.020100000e-08 V_hig
+ 5.030000000e-08 V_hig
+ 5.030100000e-08 V_hig
+ 5.040000000e-08 V_hig
+ 5.040100000e-08 V_hig
+ 5.050000000e-08 V_hig
+ 5.050100000e-08 V_hig
+ 5.060000000e-08 V_hig
+ 5.060100000e-08 V_hig
+ 5.070000000e-08 V_hig
+ 5.070100000e-08 V_hig
+ 5.080000000e-08 V_hig
+ 5.080100000e-08 V_hig
+ 5.090000000e-08 V_hig
+ 5.090100000e-08 V_low
+ 5.100000000e-08 V_low
+ 5.100100000e-08 V_low
+ 5.110000000e-08 V_low
+ 5.110100000e-08 V_low
+ 5.120000000e-08 V_low
+ 5.120100000e-08 V_low
+ 5.130000000e-08 V_low
+ 5.130100000e-08 V_low
+ 5.140000000e-08 V_low
+ 5.140100000e-08 V_low
+ 5.150000000e-08 V_low
+ 5.150100000e-08 V_low
+ 5.160000000e-08 V_low
+ 5.160100000e-08 V_low
+ 5.170000000e-08 V_low
+ 5.170100000e-08 V_low
+ 5.180000000e-08 V_low
+ 5.180100000e-08 V_low
+ 5.190000000e-08 V_low
+ 5.190100000e-08 V_low
+ 5.200000000e-08 V_low
+ 5.200100000e-08 V_low
+ 5.210000000e-08 V_low
+ 5.210100000e-08 V_low
+ 5.220000000e-08 V_low
+ 5.220100000e-08 V_low
+ 5.230000000e-08 V_low
+ 5.230100000e-08 V_low
+ 5.240000000e-08 V_low
+ 5.240100000e-08 V_low
+ 5.250000000e-08 V_low
+ 5.250100000e-08 V_low
+ 5.260000000e-08 V_low
+ 5.260100000e-08 V_low
+ 5.270000000e-08 V_low
+ 5.270100000e-08 V_low
+ 5.280000000e-08 V_low
+ 5.280100000e-08 V_low
+ 5.290000000e-08 V_low
+ 5.290100000e-08 V_hig
+ 5.300000000e-08 V_hig
+ 5.300100000e-08 V_hig
+ 5.310000000e-08 V_hig
+ 5.310100000e-08 V_hig
+ 5.320000000e-08 V_hig
+ 5.320100000e-08 V_hig
+ 5.330000000e-08 V_hig
+ 5.330100000e-08 V_hig
+ 5.340000000e-08 V_hig
+ 5.340100000e-08 V_hig
+ 5.350000000e-08 V_hig
+ 5.350100000e-08 V_hig
+ 5.360000000e-08 V_hig
+ 5.360100000e-08 V_hig
+ 5.370000000e-08 V_hig
+ 5.370100000e-08 V_hig
+ 5.380000000e-08 V_hig
+ 5.380100000e-08 V_hig
+ 5.390000000e-08 V_hig
+ 5.390100000e-08 V_low
+ 5.400000000e-08 V_low
+ 5.400100000e-08 V_low
+ 5.410000000e-08 V_low
+ 5.410100000e-08 V_low
+ 5.420000000e-08 V_low
+ 5.420100000e-08 V_low
+ 5.430000000e-08 V_low
+ 5.430100000e-08 V_low
+ 5.440000000e-08 V_low
+ 5.440100000e-08 V_low
+ 5.450000000e-08 V_low
+ 5.450100000e-08 V_low
+ 5.460000000e-08 V_low
+ 5.460100000e-08 V_low
+ 5.470000000e-08 V_low
+ 5.470100000e-08 V_low
+ 5.480000000e-08 V_low
+ 5.480100000e-08 V_low
+ 5.490000000e-08 V_low
+ 5.490100000e-08 V_hig
+ 5.500000000e-08 V_hig
+ 5.500100000e-08 V_hig
+ 5.510000000e-08 V_hig
+ 5.510100000e-08 V_hig
+ 5.520000000e-08 V_hig
+ 5.520100000e-08 V_hig
+ 5.530000000e-08 V_hig
+ 5.530100000e-08 V_hig
+ 5.540000000e-08 V_hig
+ 5.540100000e-08 V_hig
+ 5.550000000e-08 V_hig
+ 5.550100000e-08 V_hig
+ 5.560000000e-08 V_hig
+ 5.560100000e-08 V_hig
+ 5.570000000e-08 V_hig
+ 5.570100000e-08 V_hig
+ 5.580000000e-08 V_hig
+ 5.580100000e-08 V_hig
+ 5.590000000e-08 V_hig
+ 5.590100000e-08 V_hig
+ 5.600000000e-08 V_hig
+ 5.600100000e-08 V_hig
+ 5.610000000e-08 V_hig
+ 5.610100000e-08 V_hig
+ 5.620000000e-08 V_hig
+ 5.620100000e-08 V_hig
+ 5.630000000e-08 V_hig
+ 5.630100000e-08 V_hig
+ 5.640000000e-08 V_hig
+ 5.640100000e-08 V_hig
+ 5.650000000e-08 V_hig
+ 5.650100000e-08 V_hig
+ 5.660000000e-08 V_hig
+ 5.660100000e-08 V_hig
+ 5.670000000e-08 V_hig
+ 5.670100000e-08 V_hig
+ 5.680000000e-08 V_hig
+ 5.680100000e-08 V_hig
+ 5.690000000e-08 V_hig
+ 5.690100000e-08 V_hig
+ 5.700000000e-08 V_hig
+ 5.700100000e-08 V_hig
+ 5.710000000e-08 V_hig
+ 5.710100000e-08 V_hig
+ 5.720000000e-08 V_hig
+ 5.720100000e-08 V_hig
+ 5.730000000e-08 V_hig
+ 5.730100000e-08 V_hig
+ 5.740000000e-08 V_hig
+ 5.740100000e-08 V_hig
+ 5.750000000e-08 V_hig
+ 5.750100000e-08 V_hig
+ 5.760000000e-08 V_hig
+ 5.760100000e-08 V_hig
+ 5.770000000e-08 V_hig
+ 5.770100000e-08 V_hig
+ 5.780000000e-08 V_hig
+ 5.780100000e-08 V_hig
+ 5.790000000e-08 V_hig
+ 5.790100000e-08 V_hig
+ 5.800000000e-08 V_hig
+ 5.800100000e-08 V_hig
+ 5.810000000e-08 V_hig
+ 5.810100000e-08 V_hig
+ 5.820000000e-08 V_hig
+ 5.820100000e-08 V_hig
+ 5.830000000e-08 V_hig
+ 5.830100000e-08 V_hig
+ 5.840000000e-08 V_hig
+ 5.840100000e-08 V_hig
+ 5.850000000e-08 V_hig
+ 5.850100000e-08 V_hig
+ 5.860000000e-08 V_hig
+ 5.860100000e-08 V_hig
+ 5.870000000e-08 V_hig
+ 5.870100000e-08 V_hig
+ 5.880000000e-08 V_hig
+ 5.880100000e-08 V_hig
+ 5.890000000e-08 V_hig
+ 5.890100000e-08 V_low
+ 5.900000000e-08 V_low
+ 5.900100000e-08 V_low
+ 5.910000000e-08 V_low
+ 5.910100000e-08 V_low
+ 5.920000000e-08 V_low
+ 5.920100000e-08 V_low
+ 5.930000000e-08 V_low
+ 5.930100000e-08 V_low
+ 5.940000000e-08 V_low
+ 5.940100000e-08 V_low
+ 5.950000000e-08 V_low
+ 5.950100000e-08 V_low
+ 5.960000000e-08 V_low
+ 5.960100000e-08 V_low
+ 5.970000000e-08 V_low
+ 5.970100000e-08 V_low
+ 5.980000000e-08 V_low
+ 5.980100000e-08 V_low
+ 5.990000000e-08 V_low
+ 5.990100000e-08 V_low
+ 6.000000000e-08 V_low
+ 6.000100000e-08 V_low
+ 6.010000000e-08 V_low
+ 6.010100000e-08 V_low
+ 6.020000000e-08 V_low
+ 6.020100000e-08 V_low
+ 6.030000000e-08 V_low
+ 6.030100000e-08 V_low
+ 6.040000000e-08 V_low
+ 6.040100000e-08 V_low
+ 6.050000000e-08 V_low
+ 6.050100000e-08 V_low
+ 6.060000000e-08 V_low
+ 6.060100000e-08 V_low
+ 6.070000000e-08 V_low
+ 6.070100000e-08 V_low
+ 6.080000000e-08 V_low
+ 6.080100000e-08 V_low
+ 6.090000000e-08 V_low
+ 6.090100000e-08 V_hig
+ 6.100000000e-08 V_hig
+ 6.100100000e-08 V_hig
+ 6.110000000e-08 V_hig
+ 6.110100000e-08 V_hig
+ 6.120000000e-08 V_hig
+ 6.120100000e-08 V_hig
+ 6.130000000e-08 V_hig
+ 6.130100000e-08 V_hig
+ 6.140000000e-08 V_hig
+ 6.140100000e-08 V_hig
+ 6.150000000e-08 V_hig
+ 6.150100000e-08 V_hig
+ 6.160000000e-08 V_hig
+ 6.160100000e-08 V_hig
+ 6.170000000e-08 V_hig
+ 6.170100000e-08 V_hig
+ 6.180000000e-08 V_hig
+ 6.180100000e-08 V_hig
+ 6.190000000e-08 V_hig
+ 6.190100000e-08 V_hig
+ 6.200000000e-08 V_hig
+ 6.200100000e-08 V_hig
+ 6.210000000e-08 V_hig
+ 6.210100000e-08 V_hig
+ 6.220000000e-08 V_hig
+ 6.220100000e-08 V_hig
+ 6.230000000e-08 V_hig
+ 6.230100000e-08 V_hig
+ 6.240000000e-08 V_hig
+ 6.240100000e-08 V_hig
+ 6.250000000e-08 V_hig
+ 6.250100000e-08 V_hig
+ 6.260000000e-08 V_hig
+ 6.260100000e-08 V_hig
+ 6.270000000e-08 V_hig
+ 6.270100000e-08 V_hig
+ 6.280000000e-08 V_hig
+ 6.280100000e-08 V_hig
+ 6.290000000e-08 V_hig
+ 6.290100000e-08 V_low
+ 6.300000000e-08 V_low
+ 6.300100000e-08 V_low
+ 6.310000000e-08 V_low
+ 6.310100000e-08 V_low
+ 6.320000000e-08 V_low
+ 6.320100000e-08 V_low
+ 6.330000000e-08 V_low
+ 6.330100000e-08 V_low
+ 6.340000000e-08 V_low
+ 6.340100000e-08 V_low
+ 6.350000000e-08 V_low
+ 6.350100000e-08 V_low
+ 6.360000000e-08 V_low
+ 6.360100000e-08 V_low
+ 6.370000000e-08 V_low
+ 6.370100000e-08 V_low
+ 6.380000000e-08 V_low
+ 6.380100000e-08 V_low
+ 6.390000000e-08 V_low
+ 6.390100000e-08 V_low
+ 6.400000000e-08 V_low
+ 6.400100000e-08 V_low
+ 6.410000000e-08 V_low
+ 6.410100000e-08 V_low
+ 6.420000000e-08 V_low
+ 6.420100000e-08 V_low
+ 6.430000000e-08 V_low
+ 6.430100000e-08 V_low
+ 6.440000000e-08 V_low
+ 6.440100000e-08 V_low
+ 6.450000000e-08 V_low
+ 6.450100000e-08 V_low
+ 6.460000000e-08 V_low
+ 6.460100000e-08 V_low
+ 6.470000000e-08 V_low
+ 6.470100000e-08 V_low
+ 6.480000000e-08 V_low
+ 6.480100000e-08 V_low
+ 6.490000000e-08 V_low
+ 6.490100000e-08 V_hig
+ 6.500000000e-08 V_hig
+ 6.500100000e-08 V_hig
+ 6.510000000e-08 V_hig
+ 6.510100000e-08 V_hig
+ 6.520000000e-08 V_hig
+ 6.520100000e-08 V_hig
+ 6.530000000e-08 V_hig
+ 6.530100000e-08 V_hig
+ 6.540000000e-08 V_hig
+ 6.540100000e-08 V_hig
+ 6.550000000e-08 V_hig
+ 6.550100000e-08 V_hig
+ 6.560000000e-08 V_hig
+ 6.560100000e-08 V_hig
+ 6.570000000e-08 V_hig
+ 6.570100000e-08 V_hig
+ 6.580000000e-08 V_hig
+ 6.580100000e-08 V_hig
+ 6.590000000e-08 V_hig
+ 6.590100000e-08 V_hig
+ 6.600000000e-08 V_hig
+ 6.600100000e-08 V_hig
+ 6.610000000e-08 V_hig
+ 6.610100000e-08 V_hig
+ 6.620000000e-08 V_hig
+ 6.620100000e-08 V_hig
+ 6.630000000e-08 V_hig
+ 6.630100000e-08 V_hig
+ 6.640000000e-08 V_hig
+ 6.640100000e-08 V_hig
+ 6.650000000e-08 V_hig
+ 6.650100000e-08 V_hig
+ 6.660000000e-08 V_hig
+ 6.660100000e-08 V_hig
+ 6.670000000e-08 V_hig
+ 6.670100000e-08 V_hig
+ 6.680000000e-08 V_hig
+ 6.680100000e-08 V_hig
+ 6.690000000e-08 V_hig
+ 6.690100000e-08 V_low
+ 6.700000000e-08 V_low
+ 6.700100000e-08 V_low
+ 6.710000000e-08 V_low
+ 6.710100000e-08 V_low
+ 6.720000000e-08 V_low
+ 6.720100000e-08 V_low
+ 6.730000000e-08 V_low
+ 6.730100000e-08 V_low
+ 6.740000000e-08 V_low
+ 6.740100000e-08 V_low
+ 6.750000000e-08 V_low
+ 6.750100000e-08 V_low
+ 6.760000000e-08 V_low
+ 6.760100000e-08 V_low
+ 6.770000000e-08 V_low
+ 6.770100000e-08 V_low
+ 6.780000000e-08 V_low
+ 6.780100000e-08 V_low
+ 6.790000000e-08 V_low
+ 6.790100000e-08 V_low
+ 6.800000000e-08 V_low
+ 6.800100000e-08 V_low
+ 6.810000000e-08 V_low
+ 6.810100000e-08 V_low
+ 6.820000000e-08 V_low
+ 6.820100000e-08 V_low
+ 6.830000000e-08 V_low
+ 6.830100000e-08 V_low
+ 6.840000000e-08 V_low
+ 6.840100000e-08 V_low
+ 6.850000000e-08 V_low
+ 6.850100000e-08 V_low
+ 6.860000000e-08 V_low
+ 6.860100000e-08 V_low
+ 6.870000000e-08 V_low
+ 6.870100000e-08 V_low
+ 6.880000000e-08 V_low
+ 6.880100000e-08 V_low
+ 6.890000000e-08 V_low
+ 6.890100000e-08 V_low
+ 6.900000000e-08 V_low
+ 6.900100000e-08 V_low
+ 6.910000000e-08 V_low
+ 6.910100000e-08 V_low
+ 6.920000000e-08 V_low
+ 6.920100000e-08 V_low
+ 6.930000000e-08 V_low
+ 6.930100000e-08 V_low
+ 6.940000000e-08 V_low
+ 6.940100000e-08 V_low
+ 6.950000000e-08 V_low
+ 6.950100000e-08 V_low
+ 6.960000000e-08 V_low
+ 6.960100000e-08 V_low
+ 6.970000000e-08 V_low
+ 6.970100000e-08 V_low
+ 6.980000000e-08 V_low
+ 6.980100000e-08 V_low
+ 6.990000000e-08 V_low
+ 6.990100000e-08 V_hig
+ 7.000000000e-08 V_hig
+ 7.000100000e-08 V_hig
+ 7.010000000e-08 V_hig
+ 7.010100000e-08 V_hig
+ 7.020000000e-08 V_hig
+ 7.020100000e-08 V_hig
+ 7.030000000e-08 V_hig
+ 7.030100000e-08 V_hig
+ 7.040000000e-08 V_hig
+ 7.040100000e-08 V_hig
+ 7.050000000e-08 V_hig
+ 7.050100000e-08 V_hig
+ 7.060000000e-08 V_hig
+ 7.060100000e-08 V_hig
+ 7.070000000e-08 V_hig
+ 7.070100000e-08 V_hig
+ 7.080000000e-08 V_hig
+ 7.080100000e-08 V_hig
+ 7.090000000e-08 V_hig
+ 7.090100000e-08 V_low
+ 7.100000000e-08 V_low
+ 7.100100000e-08 V_low
+ 7.110000000e-08 V_low
+ 7.110100000e-08 V_low
+ 7.120000000e-08 V_low
+ 7.120100000e-08 V_low
+ 7.130000000e-08 V_low
+ 7.130100000e-08 V_low
+ 7.140000000e-08 V_low
+ 7.140100000e-08 V_low
+ 7.150000000e-08 V_low
+ 7.150100000e-08 V_low
+ 7.160000000e-08 V_low
+ 7.160100000e-08 V_low
+ 7.170000000e-08 V_low
+ 7.170100000e-08 V_low
+ 7.180000000e-08 V_low
+ 7.180100000e-08 V_low
+ 7.190000000e-08 V_low
+ 7.190100000e-08 V_hig
+ 7.200000000e-08 V_hig
+ 7.200100000e-08 V_hig
+ 7.210000000e-08 V_hig
+ 7.210100000e-08 V_hig
+ 7.220000000e-08 V_hig
+ 7.220100000e-08 V_hig
+ 7.230000000e-08 V_hig
+ 7.230100000e-08 V_hig
+ 7.240000000e-08 V_hig
+ 7.240100000e-08 V_hig
+ 7.250000000e-08 V_hig
+ 7.250100000e-08 V_hig
+ 7.260000000e-08 V_hig
+ 7.260100000e-08 V_hig
+ 7.270000000e-08 V_hig
+ 7.270100000e-08 V_hig
+ 7.280000000e-08 V_hig
+ 7.280100000e-08 V_hig
+ 7.290000000e-08 V_hig
+ 7.290100000e-08 V_low
+ 7.300000000e-08 V_low
+ 7.300100000e-08 V_low
+ 7.310000000e-08 V_low
+ 7.310100000e-08 V_low
+ 7.320000000e-08 V_low
+ 7.320100000e-08 V_low
+ 7.330000000e-08 V_low
+ 7.330100000e-08 V_low
+ 7.340000000e-08 V_low
+ 7.340100000e-08 V_low
+ 7.350000000e-08 V_low
+ 7.350100000e-08 V_low
+ 7.360000000e-08 V_low
+ 7.360100000e-08 V_low
+ 7.370000000e-08 V_low
+ 7.370100000e-08 V_low
+ 7.380000000e-08 V_low
+ 7.380100000e-08 V_low
+ 7.390000000e-08 V_low
+ 7.390100000e-08 V_hig
+ 7.400000000e-08 V_hig
+ 7.400100000e-08 V_hig
+ 7.410000000e-08 V_hig
+ 7.410100000e-08 V_hig
+ 7.420000000e-08 V_hig
+ 7.420100000e-08 V_hig
+ 7.430000000e-08 V_hig
+ 7.430100000e-08 V_hig
+ 7.440000000e-08 V_hig
+ 7.440100000e-08 V_hig
+ 7.450000000e-08 V_hig
+ 7.450100000e-08 V_hig
+ 7.460000000e-08 V_hig
+ 7.460100000e-08 V_hig
+ 7.470000000e-08 V_hig
+ 7.470100000e-08 V_hig
+ 7.480000000e-08 V_hig
+ 7.480100000e-08 V_hig
+ 7.490000000e-08 V_hig
+ 7.490100000e-08 V_low
+ 7.500000000e-08 V_low
+ 7.500100000e-08 V_low
+ 7.510000000e-08 V_low
+ 7.510100000e-08 V_low
+ 7.520000000e-08 V_low
+ 7.520100000e-08 V_low
+ 7.530000000e-08 V_low
+ 7.530100000e-08 V_low
+ 7.540000000e-08 V_low
+ 7.540100000e-08 V_low
+ 7.550000000e-08 V_low
+ 7.550100000e-08 V_low
+ 7.560000000e-08 V_low
+ 7.560100000e-08 V_low
+ 7.570000000e-08 V_low
+ 7.570100000e-08 V_low
+ 7.580000000e-08 V_low
+ 7.580100000e-08 V_low
+ 7.590000000e-08 V_low
+ 7.590100000e-08 V_low
+ 7.600000000e-08 V_low
+ 7.600100000e-08 V_low
+ 7.610000000e-08 V_low
+ 7.610100000e-08 V_low
+ 7.620000000e-08 V_low
+ 7.620100000e-08 V_low
+ 7.630000000e-08 V_low
+ 7.630100000e-08 V_low
+ 7.640000000e-08 V_low
+ 7.640100000e-08 V_low
+ 7.650000000e-08 V_low
+ 7.650100000e-08 V_low
+ 7.660000000e-08 V_low
+ 7.660100000e-08 V_low
+ 7.670000000e-08 V_low
+ 7.670100000e-08 V_low
+ 7.680000000e-08 V_low
+ 7.680100000e-08 V_low
+ 7.690000000e-08 V_low
+ 7.690100000e-08 V_hig
+ 7.700000000e-08 V_hig
+ 7.700100000e-08 V_hig
+ 7.710000000e-08 V_hig
+ 7.710100000e-08 V_hig
+ 7.720000000e-08 V_hig
+ 7.720100000e-08 V_hig
+ 7.730000000e-08 V_hig
+ 7.730100000e-08 V_hig
+ 7.740000000e-08 V_hig
+ 7.740100000e-08 V_hig
+ 7.750000000e-08 V_hig
+ 7.750100000e-08 V_hig
+ 7.760000000e-08 V_hig
+ 7.760100000e-08 V_hig
+ 7.770000000e-08 V_hig
+ 7.770100000e-08 V_hig
+ 7.780000000e-08 V_hig
+ 7.780100000e-08 V_hig
+ 7.790000000e-08 V_hig
+ 7.790100000e-08 V_hig
+ 7.800000000e-08 V_hig
+ 7.800100000e-08 V_hig
+ 7.810000000e-08 V_hig
+ 7.810100000e-08 V_hig
+ 7.820000000e-08 V_hig
+ 7.820100000e-08 V_hig
+ 7.830000000e-08 V_hig
+ 7.830100000e-08 V_hig
+ 7.840000000e-08 V_hig
+ 7.840100000e-08 V_hig
+ 7.850000000e-08 V_hig
+ 7.850100000e-08 V_hig
+ 7.860000000e-08 V_hig
+ 7.860100000e-08 V_hig
+ 7.870000000e-08 V_hig
+ 7.870100000e-08 V_hig
+ 7.880000000e-08 V_hig
+ 7.880100000e-08 V_hig
+ 7.890000000e-08 V_hig
+ 7.890100000e-08 V_low
+ 7.900000000e-08 V_low
+ 7.900100000e-08 V_low
+ 7.910000000e-08 V_low
+ 7.910100000e-08 V_low
+ 7.920000000e-08 V_low
+ 7.920100000e-08 V_low
+ 7.930000000e-08 V_low
+ 7.930100000e-08 V_low
+ 7.940000000e-08 V_low
+ 7.940100000e-08 V_low
+ 7.950000000e-08 V_low
+ 7.950100000e-08 V_low
+ 7.960000000e-08 V_low
+ 7.960100000e-08 V_low
+ 7.970000000e-08 V_low
+ 7.970100000e-08 V_low
+ 7.980000000e-08 V_low
+ 7.980100000e-08 V_low
+ 7.990000000e-08 V_low
+ 7.990100000e-08 V_low
+ 8.000000000e-08 V_low
+ 8.000100000e-08 V_low
+ 8.010000000e-08 V_low
+ 8.010100000e-08 V_low
+ 8.020000000e-08 V_low
+ 8.020100000e-08 V_low
+ 8.030000000e-08 V_low
+ 8.030100000e-08 V_low
+ 8.040000000e-08 V_low
+ 8.040100000e-08 V_low
+ 8.050000000e-08 V_low
+ 8.050100000e-08 V_low
+ 8.060000000e-08 V_low
+ 8.060100000e-08 V_low
+ 8.070000000e-08 V_low
+ 8.070100000e-08 V_low
+ 8.080000000e-08 V_low
+ 8.080100000e-08 V_low
+ 8.090000000e-08 V_low
+ 8.090100000e-08 V_hig
+ 8.100000000e-08 V_hig
+ 8.100100000e-08 V_hig
+ 8.110000000e-08 V_hig
+ 8.110100000e-08 V_hig
+ 8.120000000e-08 V_hig
+ 8.120100000e-08 V_hig
+ 8.130000000e-08 V_hig
+ 8.130100000e-08 V_hig
+ 8.140000000e-08 V_hig
+ 8.140100000e-08 V_hig
+ 8.150000000e-08 V_hig
+ 8.150100000e-08 V_hig
+ 8.160000000e-08 V_hig
+ 8.160100000e-08 V_hig
+ 8.170000000e-08 V_hig
+ 8.170100000e-08 V_hig
+ 8.180000000e-08 V_hig
+ 8.180100000e-08 V_hig
+ 8.190000000e-08 V_hig
+ 8.190100000e-08 V_hig
+ 8.200000000e-08 V_hig
+ 8.200100000e-08 V_hig
+ 8.210000000e-08 V_hig
+ 8.210100000e-08 V_hig
+ 8.220000000e-08 V_hig
+ 8.220100000e-08 V_hig
+ 8.230000000e-08 V_hig
+ 8.230100000e-08 V_hig
+ 8.240000000e-08 V_hig
+ 8.240100000e-08 V_hig
+ 8.250000000e-08 V_hig
+ 8.250100000e-08 V_hig
+ 8.260000000e-08 V_hig
+ 8.260100000e-08 V_hig
+ 8.270000000e-08 V_hig
+ 8.270100000e-08 V_hig
+ 8.280000000e-08 V_hig
+ 8.280100000e-08 V_hig
+ 8.290000000e-08 V_hig
+ 8.290100000e-08 V_low
+ 8.300000000e-08 V_low
+ 8.300100000e-08 V_low
+ 8.310000000e-08 V_low
+ 8.310100000e-08 V_low
+ 8.320000000e-08 V_low
+ 8.320100000e-08 V_low
+ 8.330000000e-08 V_low
+ 8.330100000e-08 V_low
+ 8.340000000e-08 V_low
+ 8.340100000e-08 V_low
+ 8.350000000e-08 V_low
+ 8.350100000e-08 V_low
+ 8.360000000e-08 V_low
+ 8.360100000e-08 V_low
+ 8.370000000e-08 V_low
+ 8.370100000e-08 V_low
+ 8.380000000e-08 V_low
+ 8.380100000e-08 V_low
+ 8.390000000e-08 V_low
+ 8.390100000e-08 V_low
+ 8.400000000e-08 V_low
+ 8.400100000e-08 V_low
+ 8.410000000e-08 V_low
+ 8.410100000e-08 V_low
+ 8.420000000e-08 V_low
+ 8.420100000e-08 V_low
+ 8.430000000e-08 V_low
+ 8.430100000e-08 V_low
+ 8.440000000e-08 V_low
+ 8.440100000e-08 V_low
+ 8.450000000e-08 V_low
+ 8.450100000e-08 V_low
+ 8.460000000e-08 V_low
+ 8.460100000e-08 V_low
+ 8.470000000e-08 V_low
+ 8.470100000e-08 V_low
+ 8.480000000e-08 V_low
+ 8.480100000e-08 V_low
+ 8.490000000e-08 V_low
+ 8.490100000e-08 V_low
+ 8.500000000e-08 V_low
+ 8.500100000e-08 V_low
+ 8.510000000e-08 V_low
+ 8.510100000e-08 V_low
+ 8.520000000e-08 V_low
+ 8.520100000e-08 V_low
+ 8.530000000e-08 V_low
+ 8.530100000e-08 V_low
+ 8.540000000e-08 V_low
+ 8.540100000e-08 V_low
+ 8.550000000e-08 V_low
+ 8.550100000e-08 V_low
+ 8.560000000e-08 V_low
+ 8.560100000e-08 V_low
+ 8.570000000e-08 V_low
+ 8.570100000e-08 V_low
+ 8.580000000e-08 V_low
+ 8.580100000e-08 V_low
+ 8.590000000e-08 V_low
+ 8.590100000e-08 V_low
+ 8.600000000e-08 V_low
+ 8.600100000e-08 V_low
+ 8.610000000e-08 V_low
+ 8.610100000e-08 V_low
+ 8.620000000e-08 V_low
+ 8.620100000e-08 V_low
+ 8.630000000e-08 V_low
+ 8.630100000e-08 V_low
+ 8.640000000e-08 V_low
+ 8.640100000e-08 V_low
+ 8.650000000e-08 V_low
+ 8.650100000e-08 V_low
+ 8.660000000e-08 V_low
+ 8.660100000e-08 V_low
+ 8.670000000e-08 V_low
+ 8.670100000e-08 V_low
+ 8.680000000e-08 V_low
+ 8.680100000e-08 V_low
+ 8.690000000e-08 V_low
+ 8.690100000e-08 V_hig
+ 8.700000000e-08 V_hig
+ 8.700100000e-08 V_hig
+ 8.710000000e-08 V_hig
+ 8.710100000e-08 V_hig
+ 8.720000000e-08 V_hig
+ 8.720100000e-08 V_hig
+ 8.730000000e-08 V_hig
+ 8.730100000e-08 V_hig
+ 8.740000000e-08 V_hig
+ 8.740100000e-08 V_hig
+ 8.750000000e-08 V_hig
+ 8.750100000e-08 V_hig
+ 8.760000000e-08 V_hig
+ 8.760100000e-08 V_hig
+ 8.770000000e-08 V_hig
+ 8.770100000e-08 V_hig
+ 8.780000000e-08 V_hig
+ 8.780100000e-08 V_hig
+ 8.790000000e-08 V_hig
+ 8.790100000e-08 V_hig
+ 8.800000000e-08 V_hig
+ 8.800100000e-08 V_hig
+ 8.810000000e-08 V_hig
+ 8.810100000e-08 V_hig
+ 8.820000000e-08 V_hig
+ 8.820100000e-08 V_hig
+ 8.830000000e-08 V_hig
+ 8.830100000e-08 V_hig
+ 8.840000000e-08 V_hig
+ 8.840100000e-08 V_hig
+ 8.850000000e-08 V_hig
+ 8.850100000e-08 V_hig
+ 8.860000000e-08 V_hig
+ 8.860100000e-08 V_hig
+ 8.870000000e-08 V_hig
+ 8.870100000e-08 V_hig
+ 8.880000000e-08 V_hig
+ 8.880100000e-08 V_hig
+ 8.890000000e-08 V_hig
+ 8.890100000e-08 V_hig
+ 8.900000000e-08 V_hig
+ 8.900100000e-08 V_hig
+ 8.910000000e-08 V_hig
+ 8.910100000e-08 V_hig
+ 8.920000000e-08 V_hig
+ 8.920100000e-08 V_hig
+ 8.930000000e-08 V_hig
+ 8.930100000e-08 V_hig
+ 8.940000000e-08 V_hig
+ 8.940100000e-08 V_hig
+ 8.950000000e-08 V_hig
+ 8.950100000e-08 V_hig
+ 8.960000000e-08 V_hig
+ 8.960100000e-08 V_hig
+ 8.970000000e-08 V_hig
+ 8.970100000e-08 V_hig
+ 8.980000000e-08 V_hig
+ 8.980100000e-08 V_hig
+ 8.990000000e-08 V_hig
+ 8.990100000e-08 V_low
+ 9.000000000e-08 V_low
+ 9.000100000e-08 V_low
+ 9.010000000e-08 V_low
+ 9.010100000e-08 V_low
+ 9.020000000e-08 V_low
+ 9.020100000e-08 V_low
+ 9.030000000e-08 V_low
+ 9.030100000e-08 V_low
+ 9.040000000e-08 V_low
+ 9.040100000e-08 V_low
+ 9.050000000e-08 V_low
+ 9.050100000e-08 V_low
+ 9.060000000e-08 V_low
+ 9.060100000e-08 V_low
+ 9.070000000e-08 V_low
+ 9.070100000e-08 V_low
+ 9.080000000e-08 V_low
+ 9.080100000e-08 V_low
+ 9.090000000e-08 V_low
+ 9.090100000e-08 V_low
+ 9.100000000e-08 V_low
+ 9.100100000e-08 V_low
+ 9.110000000e-08 V_low
+ 9.110100000e-08 V_low
+ 9.120000000e-08 V_low
+ 9.120100000e-08 V_low
+ 9.130000000e-08 V_low
+ 9.130100000e-08 V_low
+ 9.140000000e-08 V_low
+ 9.140100000e-08 V_low
+ 9.150000000e-08 V_low
+ 9.150100000e-08 V_low
+ 9.160000000e-08 V_low
+ 9.160100000e-08 V_low
+ 9.170000000e-08 V_low
+ 9.170100000e-08 V_low
+ 9.180000000e-08 V_low
+ 9.180100000e-08 V_low
+ 9.190000000e-08 V_low
+ 9.190100000e-08 V_low
+ 9.200000000e-08 V_low
+ 9.200100000e-08 V_low
+ 9.210000000e-08 V_low
+ 9.210100000e-08 V_low
+ 9.220000000e-08 V_low
+ 9.220100000e-08 V_low
+ 9.230000000e-08 V_low
+ 9.230100000e-08 V_low
+ 9.240000000e-08 V_low
+ 9.240100000e-08 V_low
+ 9.250000000e-08 V_low
+ 9.250100000e-08 V_low
+ 9.260000000e-08 V_low
+ 9.260100000e-08 V_low
+ 9.270000000e-08 V_low
+ 9.270100000e-08 V_low
+ 9.280000000e-08 V_low
+ 9.280100000e-08 V_low
+ 9.290000000e-08 V_low
+ 9.290100000e-08 V_hig
+ 9.300000000e-08 V_hig
+ 9.300100000e-08 V_hig
+ 9.310000000e-08 V_hig
+ 9.310100000e-08 V_hig
+ 9.320000000e-08 V_hig
+ 9.320100000e-08 V_hig
+ 9.330000000e-08 V_hig
+ 9.330100000e-08 V_hig
+ 9.340000000e-08 V_hig
+ 9.340100000e-08 V_hig
+ 9.350000000e-08 V_hig
+ 9.350100000e-08 V_hig
+ 9.360000000e-08 V_hig
+ 9.360100000e-08 V_hig
+ 9.370000000e-08 V_hig
+ 9.370100000e-08 V_hig
+ 9.380000000e-08 V_hig
+ 9.380100000e-08 V_hig
+ 9.390000000e-08 V_hig
+ 9.390100000e-08 V_hig
+ 9.400000000e-08 V_hig
+ 9.400100000e-08 V_hig
+ 9.410000000e-08 V_hig
+ 9.410100000e-08 V_hig
+ 9.420000000e-08 V_hig
+ 9.420100000e-08 V_hig
+ 9.430000000e-08 V_hig
+ 9.430100000e-08 V_hig
+ 9.440000000e-08 V_hig
+ 9.440100000e-08 V_hig
+ 9.450000000e-08 V_hig
+ 9.450100000e-08 V_hig
+ 9.460000000e-08 V_hig
+ 9.460100000e-08 V_hig
+ 9.470000000e-08 V_hig
+ 9.470100000e-08 V_hig
+ 9.480000000e-08 V_hig
+ 9.480100000e-08 V_hig
+ 9.490000000e-08 V_hig
+ 9.490100000e-08 V_hig
+ 9.500000000e-08 V_hig
+ 9.500100000e-08 V_hig
+ 9.510000000e-08 V_hig
+ 9.510100000e-08 V_hig
+ 9.520000000e-08 V_hig
+ 9.520100000e-08 V_hig
+ 9.530000000e-08 V_hig
+ 9.530100000e-08 V_hig
+ 9.540000000e-08 V_hig
+ 9.540100000e-08 V_hig
+ 9.550000000e-08 V_hig
+ 9.550100000e-08 V_hig
+ 9.560000000e-08 V_hig
+ 9.560100000e-08 V_hig
+ 9.570000000e-08 V_hig
+ 9.570100000e-08 V_hig
+ 9.580000000e-08 V_hig
+ 9.580100000e-08 V_hig
+ 9.590000000e-08 V_hig
+ 9.590100000e-08 V_low
+ 9.600000000e-08 V_low
+ 9.600100000e-08 V_low
+ 9.610000000e-08 V_low
+ 9.610100000e-08 V_low
+ 9.620000000e-08 V_low
+ 9.620100000e-08 V_low
+ 9.630000000e-08 V_low
+ 9.630100000e-08 V_low
+ 9.640000000e-08 V_low
+ 9.640100000e-08 V_low
+ 9.650000000e-08 V_low
+ 9.650100000e-08 V_low
+ 9.660000000e-08 V_low
+ 9.660100000e-08 V_low
+ 9.670000000e-08 V_low
+ 9.670100000e-08 V_low
+ 9.680000000e-08 V_low
+ 9.680100000e-08 V_low
+ 9.690000000e-08 V_low
+ 9.690100000e-08 V_low
+ 9.700000000e-08 V_low
+ 9.700100000e-08 V_low
+ 9.710000000e-08 V_low
+ 9.710100000e-08 V_low
+ 9.720000000e-08 V_low
+ 9.720100000e-08 V_low
+ 9.730000000e-08 V_low
+ 9.730100000e-08 V_low
+ 9.740000000e-08 V_low
+ 9.740100000e-08 V_low
+ 9.750000000e-08 V_low
+ 9.750100000e-08 V_low
+ 9.760000000e-08 V_low
+ 9.760100000e-08 V_low
+ 9.770000000e-08 V_low
+ 9.770100000e-08 V_low
+ 9.780000000e-08 V_low
+ 9.780100000e-08 V_low
+ 9.790000000e-08 V_low
+ 9.790100000e-08 V_low
+ 9.800000000e-08 V_low
+ 9.800100000e-08 V_low
+ 9.810000000e-08 V_low
+ 9.810100000e-08 V_low
+ 9.820000000e-08 V_low
+ 9.820100000e-08 V_low
+ 9.830000000e-08 V_low
+ 9.830100000e-08 V_low
+ 9.840000000e-08 V_low
+ 9.840100000e-08 V_low
+ 9.850000000e-08 V_low
+ 9.850100000e-08 V_low
+ 9.860000000e-08 V_low
+ 9.860100000e-08 V_low
+ 9.870000000e-08 V_low
+ 9.870100000e-08 V_low
+ 9.880000000e-08 V_low
+ 9.880100000e-08 V_low
+ 9.890000000e-08 V_low
+ 9.890100000e-08 V_low
+ 9.900000000e-08 V_low
+ 9.900100000e-08 V_low
+ 9.910000000e-08 V_low
+ 9.910100000e-08 V_low
+ 9.920000000e-08 V_low
+ 9.920100000e-08 V_low
+ 9.930000000e-08 V_low
+ 9.930100000e-08 V_low
+ 9.940000000e-08 V_low
+ 9.940100000e-08 V_low
+ 9.950000000e-08 V_low
+ 9.950100000e-08 V_low
+ 9.960000000e-08 V_low
+ 9.960100000e-08 V_low
+ 9.970000000e-08 V_low
+ 9.970100000e-08 V_low
+ 9.980000000e-08 V_low
+ 9.980100000e-08 V_low
+ 9.990000000e-08 V_low
+ 9.990100000e-08 V_hig
+ 1.000000000e-07 V_hig
+ 1.000010000e-07 V_hig
+ 1.001000000e-07 V_hig
+ 1.001010000e-07 V_hig
+ 1.002000000e-07 V_hig
+ 1.002010000e-07 V_hig
+ 1.003000000e-07 V_hig
+ 1.003010000e-07 V_hig
+ 1.004000000e-07 V_hig
+ 1.004010000e-07 V_hig
+ 1.005000000e-07 V_hig
+ 1.005010000e-07 V_hig
+ 1.006000000e-07 V_hig
+ 1.006010000e-07 V_hig
+ 1.007000000e-07 V_hig
+ 1.007010000e-07 V_hig
+ 1.008000000e-07 V_hig
+ 1.008010000e-07 V_hig
+ 1.009000000e-07 V_hig
+ 1.009010000e-07 V_low
+ 1.010000000e-07 V_low
+ 1.010010000e-07 V_low
+ 1.011000000e-07 V_low
+ 1.011010000e-07 V_low
+ 1.012000000e-07 V_low
+ 1.012010000e-07 V_low
+ 1.013000000e-07 V_low
+ 1.013010000e-07 V_low
+ 1.014000000e-07 V_low
+ 1.014010000e-07 V_low
+ 1.015000000e-07 V_low
+ 1.015010000e-07 V_low
+ 1.016000000e-07 V_low
+ 1.016010000e-07 V_low
+ 1.017000000e-07 V_low
+ 1.017010000e-07 V_low
+ 1.018000000e-07 V_low
+ 1.018010000e-07 V_low
+ 1.019000000e-07 V_low
+ 1.019010000e-07 V_hig
+ 1.020000000e-07 V_hig
+ 1.020010000e-07 V_hig
+ 1.021000000e-07 V_hig
+ 1.021010000e-07 V_hig
+ 1.022000000e-07 V_hig
+ 1.022010000e-07 V_hig
+ 1.023000000e-07 V_hig
+ 1.023010000e-07 V_hig
+ 1.024000000e-07 V_hig
+ 1.024010000e-07 V_hig
+ 1.025000000e-07 V_hig
+ 1.025010000e-07 V_hig
+ 1.026000000e-07 V_hig
+ 1.026010000e-07 V_hig
+ 1.027000000e-07 V_hig
+ 1.027010000e-07 V_hig
+ 1.028000000e-07 V_hig
+ 1.028010000e-07 V_hig
+ 1.029000000e-07 V_hig
+ 1.029010000e-07 V_hig
+ 1.030000000e-07 V_hig
+ 1.030010000e-07 V_hig
+ 1.031000000e-07 V_hig
+ 1.031010000e-07 V_hig
+ 1.032000000e-07 V_hig
+ 1.032010000e-07 V_hig
+ 1.033000000e-07 V_hig
+ 1.033010000e-07 V_hig
+ 1.034000000e-07 V_hig
+ 1.034010000e-07 V_hig
+ 1.035000000e-07 V_hig
+ 1.035010000e-07 V_hig
+ 1.036000000e-07 V_hig
+ 1.036010000e-07 V_hig
+ 1.037000000e-07 V_hig
+ 1.037010000e-07 V_hig
+ 1.038000000e-07 V_hig
+ 1.038010000e-07 V_hig
+ 1.039000000e-07 V_hig
+ 1.039010000e-07 V_low
+ 1.040000000e-07 V_low
+ 1.040010000e-07 V_low
+ 1.041000000e-07 V_low
+ 1.041010000e-07 V_low
+ 1.042000000e-07 V_low
+ 1.042010000e-07 V_low
+ 1.043000000e-07 V_low
+ 1.043010000e-07 V_low
+ 1.044000000e-07 V_low
+ 1.044010000e-07 V_low
+ 1.045000000e-07 V_low
+ 1.045010000e-07 V_low
+ 1.046000000e-07 V_low
+ 1.046010000e-07 V_low
+ 1.047000000e-07 V_low
+ 1.047010000e-07 V_low
+ 1.048000000e-07 V_low
+ 1.048010000e-07 V_low
+ 1.049000000e-07 V_low
+ 1.049010000e-07 V_low
+ 1.050000000e-07 V_low
+ 1.050010000e-07 V_low
+ 1.051000000e-07 V_low
+ 1.051010000e-07 V_low
+ 1.052000000e-07 V_low
+ 1.052010000e-07 V_low
+ 1.053000000e-07 V_low
+ 1.053010000e-07 V_low
+ 1.054000000e-07 V_low
+ 1.054010000e-07 V_low
+ 1.055000000e-07 V_low
+ 1.055010000e-07 V_low
+ 1.056000000e-07 V_low
+ 1.056010000e-07 V_low
+ 1.057000000e-07 V_low
+ 1.057010000e-07 V_low
+ 1.058000000e-07 V_low
+ 1.058010000e-07 V_low
+ 1.059000000e-07 V_low
+ 1.059010000e-07 V_low
+ 1.060000000e-07 V_low
+ 1.060010000e-07 V_low
+ 1.061000000e-07 V_low
+ 1.061010000e-07 V_low
+ 1.062000000e-07 V_low
+ 1.062010000e-07 V_low
+ 1.063000000e-07 V_low
+ 1.063010000e-07 V_low
+ 1.064000000e-07 V_low
+ 1.064010000e-07 V_low
+ 1.065000000e-07 V_low
+ 1.065010000e-07 V_low
+ 1.066000000e-07 V_low
+ 1.066010000e-07 V_low
+ 1.067000000e-07 V_low
+ 1.067010000e-07 V_low
+ 1.068000000e-07 V_low
+ 1.068010000e-07 V_low
+ 1.069000000e-07 V_low
+ 1.069010000e-07 V_hig
+ 1.070000000e-07 V_hig
+ 1.070010000e-07 V_hig
+ 1.071000000e-07 V_hig
+ 1.071010000e-07 V_hig
+ 1.072000000e-07 V_hig
+ 1.072010000e-07 V_hig
+ 1.073000000e-07 V_hig
+ 1.073010000e-07 V_hig
+ 1.074000000e-07 V_hig
+ 1.074010000e-07 V_hig
+ 1.075000000e-07 V_hig
+ 1.075010000e-07 V_hig
+ 1.076000000e-07 V_hig
+ 1.076010000e-07 V_hig
+ 1.077000000e-07 V_hig
+ 1.077010000e-07 V_hig
+ 1.078000000e-07 V_hig
+ 1.078010000e-07 V_hig
+ 1.079000000e-07 V_hig
+ 1.079010000e-07 V_low
+ 1.080000000e-07 V_low
+ 1.080010000e-07 V_low
+ 1.081000000e-07 V_low
+ 1.081010000e-07 V_low
+ 1.082000000e-07 V_low
+ 1.082010000e-07 V_low
+ 1.083000000e-07 V_low
+ 1.083010000e-07 V_low
+ 1.084000000e-07 V_low
+ 1.084010000e-07 V_low
+ 1.085000000e-07 V_low
+ 1.085010000e-07 V_low
+ 1.086000000e-07 V_low
+ 1.086010000e-07 V_low
+ 1.087000000e-07 V_low
+ 1.087010000e-07 V_low
+ 1.088000000e-07 V_low
+ 1.088010000e-07 V_low
+ 1.089000000e-07 V_low
+ 1.089010000e-07 V_low
+ 1.090000000e-07 V_low
+ 1.090010000e-07 V_low
+ 1.091000000e-07 V_low
+ 1.091010000e-07 V_low
+ 1.092000000e-07 V_low
+ 1.092010000e-07 V_low
+ 1.093000000e-07 V_low
+ 1.093010000e-07 V_low
+ 1.094000000e-07 V_low
+ 1.094010000e-07 V_low
+ 1.095000000e-07 V_low
+ 1.095010000e-07 V_low
+ 1.096000000e-07 V_low
+ 1.096010000e-07 V_low
+ 1.097000000e-07 V_low
+ 1.097010000e-07 V_low
+ 1.098000000e-07 V_low
+ 1.098010000e-07 V_low
+ 1.099000000e-07 V_low
+ 1.099010000e-07 V_hig
+ 1.100000000e-07 V_hig
+ 1.100010000e-07 V_hig
+ 1.101000000e-07 V_hig
+ 1.101010000e-07 V_hig
+ 1.102000000e-07 V_hig
+ 1.102010000e-07 V_hig
+ 1.103000000e-07 V_hig
+ 1.103010000e-07 V_hig
+ 1.104000000e-07 V_hig
+ 1.104010000e-07 V_hig
+ 1.105000000e-07 V_hig
+ 1.105010000e-07 V_hig
+ 1.106000000e-07 V_hig
+ 1.106010000e-07 V_hig
+ 1.107000000e-07 V_hig
+ 1.107010000e-07 V_hig
+ 1.108000000e-07 V_hig
+ 1.108010000e-07 V_hig
+ 1.109000000e-07 V_hig
+ 1.109010000e-07 V_low
+ 1.110000000e-07 V_low
+ 1.110010000e-07 V_low
+ 1.111000000e-07 V_low
+ 1.111010000e-07 V_low
+ 1.112000000e-07 V_low
+ 1.112010000e-07 V_low
+ 1.113000000e-07 V_low
+ 1.113010000e-07 V_low
+ 1.114000000e-07 V_low
+ 1.114010000e-07 V_low
+ 1.115000000e-07 V_low
+ 1.115010000e-07 V_low
+ 1.116000000e-07 V_low
+ 1.116010000e-07 V_low
+ 1.117000000e-07 V_low
+ 1.117010000e-07 V_low
+ 1.118000000e-07 V_low
+ 1.118010000e-07 V_low
+ 1.119000000e-07 V_low
+ 1.119010000e-07 V_hig
+ 1.120000000e-07 V_hig
+ 1.120010000e-07 V_hig
+ 1.121000000e-07 V_hig
+ 1.121010000e-07 V_hig
+ 1.122000000e-07 V_hig
+ 1.122010000e-07 V_hig
+ 1.123000000e-07 V_hig
+ 1.123010000e-07 V_hig
+ 1.124000000e-07 V_hig
+ 1.124010000e-07 V_hig
+ 1.125000000e-07 V_hig
+ 1.125010000e-07 V_hig
+ 1.126000000e-07 V_hig
+ 1.126010000e-07 V_hig
+ 1.127000000e-07 V_hig
+ 1.127010000e-07 V_hig
+ 1.128000000e-07 V_hig
+ 1.128010000e-07 V_hig
+ 1.129000000e-07 V_hig
+ 1.129010000e-07 V_low
+ 1.130000000e-07 V_low
+ 1.130010000e-07 V_low
+ 1.131000000e-07 V_low
+ 1.131010000e-07 V_low
+ 1.132000000e-07 V_low
+ 1.132010000e-07 V_low
+ 1.133000000e-07 V_low
+ 1.133010000e-07 V_low
+ 1.134000000e-07 V_low
+ 1.134010000e-07 V_low
+ 1.135000000e-07 V_low
+ 1.135010000e-07 V_low
+ 1.136000000e-07 V_low
+ 1.136010000e-07 V_low
+ 1.137000000e-07 V_low
+ 1.137010000e-07 V_low
+ 1.138000000e-07 V_low
+ 1.138010000e-07 V_low
+ 1.139000000e-07 V_low
+ 1.139010000e-07 V_hig
+ 1.140000000e-07 V_hig
+ 1.140010000e-07 V_hig
+ 1.141000000e-07 V_hig
+ 1.141010000e-07 V_hig
+ 1.142000000e-07 V_hig
+ 1.142010000e-07 V_hig
+ 1.143000000e-07 V_hig
+ 1.143010000e-07 V_hig
+ 1.144000000e-07 V_hig
+ 1.144010000e-07 V_hig
+ 1.145000000e-07 V_hig
+ 1.145010000e-07 V_hig
+ 1.146000000e-07 V_hig
+ 1.146010000e-07 V_hig
+ 1.147000000e-07 V_hig
+ 1.147010000e-07 V_hig
+ 1.148000000e-07 V_hig
+ 1.148010000e-07 V_hig
+ 1.149000000e-07 V_hig
+ 1.149010000e-07 V_hig
+ 1.150000000e-07 V_hig
+ 1.150010000e-07 V_hig
+ 1.151000000e-07 V_hig
+ 1.151010000e-07 V_hig
+ 1.152000000e-07 V_hig
+ 1.152010000e-07 V_hig
+ 1.153000000e-07 V_hig
+ 1.153010000e-07 V_hig
+ 1.154000000e-07 V_hig
+ 1.154010000e-07 V_hig
+ 1.155000000e-07 V_hig
+ 1.155010000e-07 V_hig
+ 1.156000000e-07 V_hig
+ 1.156010000e-07 V_hig
+ 1.157000000e-07 V_hig
+ 1.157010000e-07 V_hig
+ 1.158000000e-07 V_hig
+ 1.158010000e-07 V_hig
+ 1.159000000e-07 V_hig
+ 1.159010000e-07 V_low
+ 1.160000000e-07 V_low
+ 1.160010000e-07 V_low
+ 1.161000000e-07 V_low
+ 1.161010000e-07 V_low
+ 1.162000000e-07 V_low
+ 1.162010000e-07 V_low
+ 1.163000000e-07 V_low
+ 1.163010000e-07 V_low
+ 1.164000000e-07 V_low
+ 1.164010000e-07 V_low
+ 1.165000000e-07 V_low
+ 1.165010000e-07 V_low
+ 1.166000000e-07 V_low
+ 1.166010000e-07 V_low
+ 1.167000000e-07 V_low
+ 1.167010000e-07 V_low
+ 1.168000000e-07 V_low
+ 1.168010000e-07 V_low
+ 1.169000000e-07 V_low
+ 1.169010000e-07 V_hig
+ 1.170000000e-07 V_hig
+ 1.170010000e-07 V_hig
+ 1.171000000e-07 V_hig
+ 1.171010000e-07 V_hig
+ 1.172000000e-07 V_hig
+ 1.172010000e-07 V_hig
+ 1.173000000e-07 V_hig
+ 1.173010000e-07 V_hig
+ 1.174000000e-07 V_hig
+ 1.174010000e-07 V_hig
+ 1.175000000e-07 V_hig
+ 1.175010000e-07 V_hig
+ 1.176000000e-07 V_hig
+ 1.176010000e-07 V_hig
+ 1.177000000e-07 V_hig
+ 1.177010000e-07 V_hig
+ 1.178000000e-07 V_hig
+ 1.178010000e-07 V_hig
+ 1.179000000e-07 V_hig
+ 1.179010000e-07 V_hig
+ 1.180000000e-07 V_hig
+ 1.180010000e-07 V_hig
+ 1.181000000e-07 V_hig
+ 1.181010000e-07 V_hig
+ 1.182000000e-07 V_hig
+ 1.182010000e-07 V_hig
+ 1.183000000e-07 V_hig
+ 1.183010000e-07 V_hig
+ 1.184000000e-07 V_hig
+ 1.184010000e-07 V_hig
+ 1.185000000e-07 V_hig
+ 1.185010000e-07 V_hig
+ 1.186000000e-07 V_hig
+ 1.186010000e-07 V_hig
+ 1.187000000e-07 V_hig
+ 1.187010000e-07 V_hig
+ 1.188000000e-07 V_hig
+ 1.188010000e-07 V_hig
+ 1.189000000e-07 V_hig
+ 1.189010000e-07 V_low
+ 1.190000000e-07 V_low
+ 1.190010000e-07 V_low
+ 1.191000000e-07 V_low
+ 1.191010000e-07 V_low
+ 1.192000000e-07 V_low
+ 1.192010000e-07 V_low
+ 1.193000000e-07 V_low
+ 1.193010000e-07 V_low
+ 1.194000000e-07 V_low
+ 1.194010000e-07 V_low
+ 1.195000000e-07 V_low
+ 1.195010000e-07 V_low
+ 1.196000000e-07 V_low
+ 1.196010000e-07 V_low
+ 1.197000000e-07 V_low
+ 1.197010000e-07 V_low
+ 1.198000000e-07 V_low
+ 1.198010000e-07 V_low
+ 1.199000000e-07 V_low
+ 1.199010000e-07 V_hig
+ 1.200000000e-07 V_hig
+ 1.200010000e-07 V_hig
+ 1.201000000e-07 V_hig
+ 1.201010000e-07 V_hig
+ 1.202000000e-07 V_hig
+ 1.202010000e-07 V_hig
+ 1.203000000e-07 V_hig
+ 1.203010000e-07 V_hig
+ 1.204000000e-07 V_hig
+ 1.204010000e-07 V_hig
+ 1.205000000e-07 V_hig
+ 1.205010000e-07 V_hig
+ 1.206000000e-07 V_hig
+ 1.206010000e-07 V_hig
+ 1.207000000e-07 V_hig
+ 1.207010000e-07 V_hig
+ 1.208000000e-07 V_hig
+ 1.208010000e-07 V_hig
+ 1.209000000e-07 V_hig
+ 1.209010000e-07 V_hig
+ 1.210000000e-07 V_hig
+ 1.210010000e-07 V_hig
+ 1.211000000e-07 V_hig
+ 1.211010000e-07 V_hig
+ 1.212000000e-07 V_hig
+ 1.212010000e-07 V_hig
+ 1.213000000e-07 V_hig
+ 1.213010000e-07 V_hig
+ 1.214000000e-07 V_hig
+ 1.214010000e-07 V_hig
+ 1.215000000e-07 V_hig
+ 1.215010000e-07 V_hig
+ 1.216000000e-07 V_hig
+ 1.216010000e-07 V_hig
+ 1.217000000e-07 V_hig
+ 1.217010000e-07 V_hig
+ 1.218000000e-07 V_hig
+ 1.218010000e-07 V_hig
+ 1.219000000e-07 V_hig
+ 1.219010000e-07 V_low
+ 1.220000000e-07 V_low
+ 1.220010000e-07 V_low
+ 1.221000000e-07 V_low
+ 1.221010000e-07 V_low
+ 1.222000000e-07 V_low
+ 1.222010000e-07 V_low
+ 1.223000000e-07 V_low
+ 1.223010000e-07 V_low
+ 1.224000000e-07 V_low
+ 1.224010000e-07 V_low
+ 1.225000000e-07 V_low
+ 1.225010000e-07 V_low
+ 1.226000000e-07 V_low
+ 1.226010000e-07 V_low
+ 1.227000000e-07 V_low
+ 1.227010000e-07 V_low
+ 1.228000000e-07 V_low
+ 1.228010000e-07 V_low
+ 1.229000000e-07 V_low
+ 1.229010000e-07 V_hig
+ 1.230000000e-07 V_hig
+ 1.230010000e-07 V_hig
+ 1.231000000e-07 V_hig
+ 1.231010000e-07 V_hig
+ 1.232000000e-07 V_hig
+ 1.232010000e-07 V_hig
+ 1.233000000e-07 V_hig
+ 1.233010000e-07 V_hig
+ 1.234000000e-07 V_hig
+ 1.234010000e-07 V_hig
+ 1.235000000e-07 V_hig
+ 1.235010000e-07 V_hig
+ 1.236000000e-07 V_hig
+ 1.236010000e-07 V_hig
+ 1.237000000e-07 V_hig
+ 1.237010000e-07 V_hig
+ 1.238000000e-07 V_hig
+ 1.238010000e-07 V_hig
+ 1.239000000e-07 V_hig
+ 1.239010000e-07 V_low
+ 1.240000000e-07 V_low
+ 1.240010000e-07 V_low
+ 1.241000000e-07 V_low
+ 1.241010000e-07 V_low
+ 1.242000000e-07 V_low
+ 1.242010000e-07 V_low
+ 1.243000000e-07 V_low
+ 1.243010000e-07 V_low
+ 1.244000000e-07 V_low
+ 1.244010000e-07 V_low
+ 1.245000000e-07 V_low
+ 1.245010000e-07 V_low
+ 1.246000000e-07 V_low
+ 1.246010000e-07 V_low
+ 1.247000000e-07 V_low
+ 1.247010000e-07 V_low
+ 1.248000000e-07 V_low
+ 1.248010000e-07 V_low
+ 1.249000000e-07 V_low
+ 1.249010000e-07 V_hig
+ 1.250000000e-07 V_hig
+ 1.250010000e-07 V_hig
+ 1.251000000e-07 V_hig
+ 1.251010000e-07 V_hig
+ 1.252000000e-07 V_hig
+ 1.252010000e-07 V_hig
+ 1.253000000e-07 V_hig
+ 1.253010000e-07 V_hig
+ 1.254000000e-07 V_hig
+ 1.254010000e-07 V_hig
+ 1.255000000e-07 V_hig
+ 1.255010000e-07 V_hig
+ 1.256000000e-07 V_hig
+ 1.256010000e-07 V_hig
+ 1.257000000e-07 V_hig
+ 1.257010000e-07 V_hig
+ 1.258000000e-07 V_hig
+ 1.258010000e-07 V_hig
+ 1.259000000e-07 V_hig
+ 1.259010000e-07 V_low
+ 1.260000000e-07 V_low
+ 1.260010000e-07 V_low
+ 1.261000000e-07 V_low
+ 1.261010000e-07 V_low
+ 1.262000000e-07 V_low
+ 1.262010000e-07 V_low
+ 1.263000000e-07 V_low
+ 1.263010000e-07 V_low
+ 1.264000000e-07 V_low
+ 1.264010000e-07 V_low
+ 1.265000000e-07 V_low
+ 1.265010000e-07 V_low
+ 1.266000000e-07 V_low
+ 1.266010000e-07 V_low
+ 1.267000000e-07 V_low
+ 1.267010000e-07 V_low
+ 1.268000000e-07 V_low
+ 1.268010000e-07 V_low
+ 1.269000000e-07 V_low
+ 1.269010000e-07 V_hig
+ 1.270000000e-07 V_hig
+ 1.270010000e-07 V_hig
+ 1.271000000e-07 V_hig
+ 1.271010000e-07 V_hig
+ 1.272000000e-07 V_hig
+ 1.272010000e-07 V_hig
+ 1.273000000e-07 V_hig
+ 1.273010000e-07 V_hig
+ 1.274000000e-07 V_hig
+ 1.274010000e-07 V_hig
+ 1.275000000e-07 V_hig
+ 1.275010000e-07 V_hig
+ 1.276000000e-07 V_hig
+ 1.276010000e-07 V_hig
+ 1.277000000e-07 V_hig
+ 1.277010000e-07 V_hig
+ 1.278000000e-07 V_hig
+ 1.278010000e-07 V_hig
+ 1.279000000e-07 V_hig
+ 1.279010000e-07 V_hig
+ 1.280000000e-07 V_hig
+ 1.280010000e-07 V_hig
+ 1.281000000e-07 V_hig
+ 1.281010000e-07 V_hig
+ 1.282000000e-07 V_hig
+ 1.282010000e-07 V_hig
+ 1.283000000e-07 V_hig
+ 1.283010000e-07 V_hig
+ 1.284000000e-07 V_hig
+ 1.284010000e-07 V_hig
+ 1.285000000e-07 V_hig
+ 1.285010000e-07 V_hig
+ 1.286000000e-07 V_hig
+ 1.286010000e-07 V_hig
+ 1.287000000e-07 V_hig
+ 1.287010000e-07 V_hig
+ 1.288000000e-07 V_hig
+ 1.288010000e-07 V_hig
+ 1.289000000e-07 V_hig
+ 1.289010000e-07 V_low
+ 1.290000000e-07 V_low
+ 1.290010000e-07 V_low
+ 1.291000000e-07 V_low
+ 1.291010000e-07 V_low
+ 1.292000000e-07 V_low
+ 1.292010000e-07 V_low
+ 1.293000000e-07 V_low
+ 1.293010000e-07 V_low
+ 1.294000000e-07 V_low
+ 1.294010000e-07 V_low
+ 1.295000000e-07 V_low
+ 1.295010000e-07 V_low
+ 1.296000000e-07 V_low
+ 1.296010000e-07 V_low
+ 1.297000000e-07 V_low
+ 1.297010000e-07 V_low
+ 1.298000000e-07 V_low
+ 1.298010000e-07 V_low
+ 1.299000000e-07 V_low
+ 1.299010000e-07 V_hig
+ 1.300000000e-07 V_hig
+ 1.300010000e-07 V_hig
+ 1.301000000e-07 V_hig
+ 1.301010000e-07 V_hig
+ 1.302000000e-07 V_hig
+ 1.302010000e-07 V_hig
+ 1.303000000e-07 V_hig
+ 1.303010000e-07 V_hig
+ 1.304000000e-07 V_hig
+ 1.304010000e-07 V_hig
+ 1.305000000e-07 V_hig
+ 1.305010000e-07 V_hig
+ 1.306000000e-07 V_hig
+ 1.306010000e-07 V_hig
+ 1.307000000e-07 V_hig
+ 1.307010000e-07 V_hig
+ 1.308000000e-07 V_hig
+ 1.308010000e-07 V_hig
+ 1.309000000e-07 V_hig
+ 1.309010000e-07 V_low
+ 1.310000000e-07 V_low
+ 1.310010000e-07 V_low
+ 1.311000000e-07 V_low
+ 1.311010000e-07 V_low
+ 1.312000000e-07 V_low
+ 1.312010000e-07 V_low
+ 1.313000000e-07 V_low
+ 1.313010000e-07 V_low
+ 1.314000000e-07 V_low
+ 1.314010000e-07 V_low
+ 1.315000000e-07 V_low
+ 1.315010000e-07 V_low
+ 1.316000000e-07 V_low
+ 1.316010000e-07 V_low
+ 1.317000000e-07 V_low
+ 1.317010000e-07 V_low
+ 1.318000000e-07 V_low
+ 1.318010000e-07 V_low
+ 1.319000000e-07 V_low
+ 1.319010000e-07 V_low
+ 1.320000000e-07 V_low
+ 1.320010000e-07 V_low
+ 1.321000000e-07 V_low
+ 1.321010000e-07 V_low
+ 1.322000000e-07 V_low
+ 1.322010000e-07 V_low
+ 1.323000000e-07 V_low
+ 1.323010000e-07 V_low
+ 1.324000000e-07 V_low
+ 1.324010000e-07 V_low
+ 1.325000000e-07 V_low
+ 1.325010000e-07 V_low
+ 1.326000000e-07 V_low
+ 1.326010000e-07 V_low
+ 1.327000000e-07 V_low
+ 1.327010000e-07 V_low
+ 1.328000000e-07 V_low
+ 1.328010000e-07 V_low
+ 1.329000000e-07 V_low
+ 1.329010000e-07 V_low
+ 1.330000000e-07 V_low
+ 1.330010000e-07 V_low
+ 1.331000000e-07 V_low
+ 1.331010000e-07 V_low
+ 1.332000000e-07 V_low
+ 1.332010000e-07 V_low
+ 1.333000000e-07 V_low
+ 1.333010000e-07 V_low
+ 1.334000000e-07 V_low
+ 1.334010000e-07 V_low
+ 1.335000000e-07 V_low
+ 1.335010000e-07 V_low
+ 1.336000000e-07 V_low
+ 1.336010000e-07 V_low
+ 1.337000000e-07 V_low
+ 1.337010000e-07 V_low
+ 1.338000000e-07 V_low
+ 1.338010000e-07 V_low
+ 1.339000000e-07 V_low
+ 1.339010000e-07 V_hig
+ 1.340000000e-07 V_hig
+ 1.340010000e-07 V_hig
+ 1.341000000e-07 V_hig
+ 1.341010000e-07 V_hig
+ 1.342000000e-07 V_hig
+ 1.342010000e-07 V_hig
+ 1.343000000e-07 V_hig
+ 1.343010000e-07 V_hig
+ 1.344000000e-07 V_hig
+ 1.344010000e-07 V_hig
+ 1.345000000e-07 V_hig
+ 1.345010000e-07 V_hig
+ 1.346000000e-07 V_hig
+ 1.346010000e-07 V_hig
+ 1.347000000e-07 V_hig
+ 1.347010000e-07 V_hig
+ 1.348000000e-07 V_hig
+ 1.348010000e-07 V_hig
+ 1.349000000e-07 V_hig
+ 1.349010000e-07 V_hig
+ 1.350000000e-07 V_hig
+ 1.350010000e-07 V_hig
+ 1.351000000e-07 V_hig
+ 1.351010000e-07 V_hig
+ 1.352000000e-07 V_hig
+ 1.352010000e-07 V_hig
+ 1.353000000e-07 V_hig
+ 1.353010000e-07 V_hig
+ 1.354000000e-07 V_hig
+ 1.354010000e-07 V_hig
+ 1.355000000e-07 V_hig
+ 1.355010000e-07 V_hig
+ 1.356000000e-07 V_hig
+ 1.356010000e-07 V_hig
+ 1.357000000e-07 V_hig
+ 1.357010000e-07 V_hig
+ 1.358000000e-07 V_hig
+ 1.358010000e-07 V_hig
+ 1.359000000e-07 V_hig
+ 1.359010000e-07 V_hig
+ 1.360000000e-07 V_hig
+ 1.360010000e-07 V_hig
+ 1.361000000e-07 V_hig
+ 1.361010000e-07 V_hig
+ 1.362000000e-07 V_hig
+ 1.362010000e-07 V_hig
+ 1.363000000e-07 V_hig
+ 1.363010000e-07 V_hig
+ 1.364000000e-07 V_hig
+ 1.364010000e-07 V_hig
+ 1.365000000e-07 V_hig
+ 1.365010000e-07 V_hig
+ 1.366000000e-07 V_hig
+ 1.366010000e-07 V_hig
+ 1.367000000e-07 V_hig
+ 1.367010000e-07 V_hig
+ 1.368000000e-07 V_hig
+ 1.368010000e-07 V_hig
+ 1.369000000e-07 V_hig
+ 1.369010000e-07 V_hig
+ 1.370000000e-07 V_hig
+ 1.370010000e-07 V_hig
+ 1.371000000e-07 V_hig
+ 1.371010000e-07 V_hig
+ 1.372000000e-07 V_hig
+ 1.372010000e-07 V_hig
+ 1.373000000e-07 V_hig
+ 1.373010000e-07 V_hig
+ 1.374000000e-07 V_hig
+ 1.374010000e-07 V_hig
+ 1.375000000e-07 V_hig
+ 1.375010000e-07 V_hig
+ 1.376000000e-07 V_hig
+ 1.376010000e-07 V_hig
+ 1.377000000e-07 V_hig
+ 1.377010000e-07 V_hig
+ 1.378000000e-07 V_hig
+ 1.378010000e-07 V_hig
+ 1.379000000e-07 V_hig
+ 1.379010000e-07 V_hig
+ 1.380000000e-07 V_hig
+ 1.380010000e-07 V_hig
+ 1.381000000e-07 V_hig
+ 1.381010000e-07 V_hig
+ 1.382000000e-07 V_hig
+ 1.382010000e-07 V_hig
+ 1.383000000e-07 V_hig
+ 1.383010000e-07 V_hig
+ 1.384000000e-07 V_hig
+ 1.384010000e-07 V_hig
+ 1.385000000e-07 V_hig
+ 1.385010000e-07 V_hig
+ 1.386000000e-07 V_hig
+ 1.386010000e-07 V_hig
+ 1.387000000e-07 V_hig
+ 1.387010000e-07 V_hig
+ 1.388000000e-07 V_hig
+ 1.388010000e-07 V_hig
+ 1.389000000e-07 V_hig
+ 1.389010000e-07 V_low
+ 1.390000000e-07 V_low
+ 1.390010000e-07 V_low
+ 1.391000000e-07 V_low
+ 1.391010000e-07 V_low
+ 1.392000000e-07 V_low
+ 1.392010000e-07 V_low
+ 1.393000000e-07 V_low
+ 1.393010000e-07 V_low
+ 1.394000000e-07 V_low
+ 1.394010000e-07 V_low
+ 1.395000000e-07 V_low
+ 1.395010000e-07 V_low
+ 1.396000000e-07 V_low
+ 1.396010000e-07 V_low
+ 1.397000000e-07 V_low
+ 1.397010000e-07 V_low
+ 1.398000000e-07 V_low
+ 1.398010000e-07 V_low
+ 1.399000000e-07 V_low
+ 1.399010000e-07 V_hig
+ 1.400000000e-07 V_hig
+ 1.400010000e-07 V_hig
+ 1.401000000e-07 V_hig
+ 1.401010000e-07 V_hig
+ 1.402000000e-07 V_hig
+ 1.402010000e-07 V_hig
+ 1.403000000e-07 V_hig
+ 1.403010000e-07 V_hig
+ 1.404000000e-07 V_hig
+ 1.404010000e-07 V_hig
+ 1.405000000e-07 V_hig
+ 1.405010000e-07 V_hig
+ 1.406000000e-07 V_hig
+ 1.406010000e-07 V_hig
+ 1.407000000e-07 V_hig
+ 1.407010000e-07 V_hig
+ 1.408000000e-07 V_hig
+ 1.408010000e-07 V_hig
+ 1.409000000e-07 V_hig
+ 1.409010000e-07 V_low
+ 1.410000000e-07 V_low
+ 1.410010000e-07 V_low
+ 1.411000000e-07 V_low
+ 1.411010000e-07 V_low
+ 1.412000000e-07 V_low
+ 1.412010000e-07 V_low
+ 1.413000000e-07 V_low
+ 1.413010000e-07 V_low
+ 1.414000000e-07 V_low
+ 1.414010000e-07 V_low
+ 1.415000000e-07 V_low
+ 1.415010000e-07 V_low
+ 1.416000000e-07 V_low
+ 1.416010000e-07 V_low
+ 1.417000000e-07 V_low
+ 1.417010000e-07 V_low
+ 1.418000000e-07 V_low
+ 1.418010000e-07 V_low
+ 1.419000000e-07 V_low
+ 1.419010000e-07 V_hig
+ 1.420000000e-07 V_hig
+ 1.420010000e-07 V_hig
+ 1.421000000e-07 V_hig
+ 1.421010000e-07 V_hig
+ 1.422000000e-07 V_hig
+ 1.422010000e-07 V_hig
+ 1.423000000e-07 V_hig
+ 1.423010000e-07 V_hig
+ 1.424000000e-07 V_hig
+ 1.424010000e-07 V_hig
+ 1.425000000e-07 V_hig
+ 1.425010000e-07 V_hig
+ 1.426000000e-07 V_hig
+ 1.426010000e-07 V_hig
+ 1.427000000e-07 V_hig
+ 1.427010000e-07 V_hig
+ 1.428000000e-07 V_hig
+ 1.428010000e-07 V_hig
+ 1.429000000e-07 V_hig
+ 1.429010000e-07 V_low
+ 1.430000000e-07 V_low
+ 1.430010000e-07 V_low
+ 1.431000000e-07 V_low
+ 1.431010000e-07 V_low
+ 1.432000000e-07 V_low
+ 1.432010000e-07 V_low
+ 1.433000000e-07 V_low
+ 1.433010000e-07 V_low
+ 1.434000000e-07 V_low
+ 1.434010000e-07 V_low
+ 1.435000000e-07 V_low
+ 1.435010000e-07 V_low
+ 1.436000000e-07 V_low
+ 1.436010000e-07 V_low
+ 1.437000000e-07 V_low
+ 1.437010000e-07 V_low
+ 1.438000000e-07 V_low
+ 1.438010000e-07 V_low
+ 1.439000000e-07 V_low
+ 1.439010000e-07 V_low
+ 1.440000000e-07 V_low
+ 1.440010000e-07 V_low
+ 1.441000000e-07 V_low
+ 1.441010000e-07 V_low
+ 1.442000000e-07 V_low
+ 1.442010000e-07 V_low
+ 1.443000000e-07 V_low
+ 1.443010000e-07 V_low
+ 1.444000000e-07 V_low
+ 1.444010000e-07 V_low
+ 1.445000000e-07 V_low
+ 1.445010000e-07 V_low
+ 1.446000000e-07 V_low
+ 1.446010000e-07 V_low
+ 1.447000000e-07 V_low
+ 1.447010000e-07 V_low
+ 1.448000000e-07 V_low
+ 1.448010000e-07 V_low
+ 1.449000000e-07 V_low
+ 1.449010000e-07 V_low
+ 1.450000000e-07 V_low
+ 1.450010000e-07 V_low
+ 1.451000000e-07 V_low
+ 1.451010000e-07 V_low
+ 1.452000000e-07 V_low
+ 1.452010000e-07 V_low
+ 1.453000000e-07 V_low
+ 1.453010000e-07 V_low
+ 1.454000000e-07 V_low
+ 1.454010000e-07 V_low
+ 1.455000000e-07 V_low
+ 1.455010000e-07 V_low
+ 1.456000000e-07 V_low
+ 1.456010000e-07 V_low
+ 1.457000000e-07 V_low
+ 1.457010000e-07 V_low
+ 1.458000000e-07 V_low
+ 1.458010000e-07 V_low
+ 1.459000000e-07 V_low
+ 1.459010000e-07 V_hig
+ 1.460000000e-07 V_hig
+ 1.460010000e-07 V_hig
+ 1.461000000e-07 V_hig
+ 1.461010000e-07 V_hig
+ 1.462000000e-07 V_hig
+ 1.462010000e-07 V_hig
+ 1.463000000e-07 V_hig
+ 1.463010000e-07 V_hig
+ 1.464000000e-07 V_hig
+ 1.464010000e-07 V_hig
+ 1.465000000e-07 V_hig
+ 1.465010000e-07 V_hig
+ 1.466000000e-07 V_hig
+ 1.466010000e-07 V_hig
+ 1.467000000e-07 V_hig
+ 1.467010000e-07 V_hig
+ 1.468000000e-07 V_hig
+ 1.468010000e-07 V_hig
+ 1.469000000e-07 V_hig
+ 1.469010000e-07 V_hig
+ 1.470000000e-07 V_hig
+ 1.470010000e-07 V_hig
+ 1.471000000e-07 V_hig
+ 1.471010000e-07 V_hig
+ 1.472000000e-07 V_hig
+ 1.472010000e-07 V_hig
+ 1.473000000e-07 V_hig
+ 1.473010000e-07 V_hig
+ 1.474000000e-07 V_hig
+ 1.474010000e-07 V_hig
+ 1.475000000e-07 V_hig
+ 1.475010000e-07 V_hig
+ 1.476000000e-07 V_hig
+ 1.476010000e-07 V_hig
+ 1.477000000e-07 V_hig
+ 1.477010000e-07 V_hig
+ 1.478000000e-07 V_hig
+ 1.478010000e-07 V_hig
+ 1.479000000e-07 V_hig
+ 1.479010000e-07 V_low
+ 1.480000000e-07 V_low
+ 1.480010000e-07 V_low
+ 1.481000000e-07 V_low
+ 1.481010000e-07 V_low
+ 1.482000000e-07 V_low
+ 1.482010000e-07 V_low
+ 1.483000000e-07 V_low
+ 1.483010000e-07 V_low
+ 1.484000000e-07 V_low
+ 1.484010000e-07 V_low
+ 1.485000000e-07 V_low
+ 1.485010000e-07 V_low
+ 1.486000000e-07 V_low
+ 1.486010000e-07 V_low
+ 1.487000000e-07 V_low
+ 1.487010000e-07 V_low
+ 1.488000000e-07 V_low
+ 1.488010000e-07 V_low
+ 1.489000000e-07 V_low
+ 1.489010000e-07 V_hig
+ 1.490000000e-07 V_hig
+ 1.490010000e-07 V_hig
+ 1.491000000e-07 V_hig
+ 1.491010000e-07 V_hig
+ 1.492000000e-07 V_hig
+ 1.492010000e-07 V_hig
+ 1.493000000e-07 V_hig
+ 1.493010000e-07 V_hig
+ 1.494000000e-07 V_hig
+ 1.494010000e-07 V_hig
+ 1.495000000e-07 V_hig
+ 1.495010000e-07 V_hig
+ 1.496000000e-07 V_hig
+ 1.496010000e-07 V_hig
+ 1.497000000e-07 V_hig
+ 1.497010000e-07 V_hig
+ 1.498000000e-07 V_hig
+ 1.498010000e-07 V_hig
+ 1.499000000e-07 V_hig
+ 1.499010000e-07 V_low
+ 1.500000000e-07 V_low
+ 1.500010000e-07 V_low
+ 1.501000000e-07 V_low
+ 1.501010000e-07 V_low
+ 1.502000000e-07 V_low
+ 1.502010000e-07 V_low
+ 1.503000000e-07 V_low
+ 1.503010000e-07 V_low
+ 1.504000000e-07 V_low
+ 1.504010000e-07 V_low
+ 1.505000000e-07 V_low
+ 1.505010000e-07 V_low
+ 1.506000000e-07 V_low
+ 1.506010000e-07 V_low
+ 1.507000000e-07 V_low
+ 1.507010000e-07 V_low
+ 1.508000000e-07 V_low
+ 1.508010000e-07 V_low
+ 1.509000000e-07 V_low
+ 1.509010000e-07 V_low
+ 1.510000000e-07 V_low
+ 1.510010000e-07 V_low
+ 1.511000000e-07 V_low
+ 1.511010000e-07 V_low
+ 1.512000000e-07 V_low
+ 1.512010000e-07 V_low
+ 1.513000000e-07 V_low
+ 1.513010000e-07 V_low
+ 1.514000000e-07 V_low
+ 1.514010000e-07 V_low
+ 1.515000000e-07 V_low
+ 1.515010000e-07 V_low
+ 1.516000000e-07 V_low
+ 1.516010000e-07 V_low
+ 1.517000000e-07 V_low
+ 1.517010000e-07 V_low
+ 1.518000000e-07 V_low
+ 1.518010000e-07 V_low
+ 1.519000000e-07 V_low
+ 1.519010000e-07 V_low
+ 1.520000000e-07 V_low
+ 1.520010000e-07 V_low
+ 1.521000000e-07 V_low
+ 1.521010000e-07 V_low
+ 1.522000000e-07 V_low
+ 1.522010000e-07 V_low
+ 1.523000000e-07 V_low
+ 1.523010000e-07 V_low
+ 1.524000000e-07 V_low
+ 1.524010000e-07 V_low
+ 1.525000000e-07 V_low
+ 1.525010000e-07 V_low
+ 1.526000000e-07 V_low
+ 1.526010000e-07 V_low
+ 1.527000000e-07 V_low
+ 1.527010000e-07 V_low
+ 1.528000000e-07 V_low
+ 1.528010000e-07 V_low
+ 1.529000000e-07 V_low
+ 1.529010000e-07 V_low
+ 1.530000000e-07 V_low
+ 1.530010000e-07 V_low
+ 1.531000000e-07 V_low
+ 1.531010000e-07 V_low
+ 1.532000000e-07 V_low
+ 1.532010000e-07 V_low
+ 1.533000000e-07 V_low
+ 1.533010000e-07 V_low
+ 1.534000000e-07 V_low
+ 1.534010000e-07 V_low
+ 1.535000000e-07 V_low
+ 1.535010000e-07 V_low
+ 1.536000000e-07 V_low
+ 1.536010000e-07 V_low
+ 1.537000000e-07 V_low
+ 1.537010000e-07 V_low
+ 1.538000000e-07 V_low
+ 1.538010000e-07 V_low
+ 1.539000000e-07 V_low
+ 1.539010000e-07 V_low
+ 1.540000000e-07 V_low
+ 1.540010000e-07 V_low
+ 1.541000000e-07 V_low
+ 1.541010000e-07 V_low
+ 1.542000000e-07 V_low
+ 1.542010000e-07 V_low
+ 1.543000000e-07 V_low
+ 1.543010000e-07 V_low
+ 1.544000000e-07 V_low
+ 1.544010000e-07 V_low
+ 1.545000000e-07 V_low
+ 1.545010000e-07 V_low
+ 1.546000000e-07 V_low
+ 1.546010000e-07 V_low
+ 1.547000000e-07 V_low
+ 1.547010000e-07 V_low
+ 1.548000000e-07 V_low
+ 1.548010000e-07 V_low
+ 1.549000000e-07 V_low
+ 1.549010000e-07 V_hig
+ 1.550000000e-07 V_hig
+ 1.550010000e-07 V_hig
+ 1.551000000e-07 V_hig
+ 1.551010000e-07 V_hig
+ 1.552000000e-07 V_hig
+ 1.552010000e-07 V_hig
+ 1.553000000e-07 V_hig
+ 1.553010000e-07 V_hig
+ 1.554000000e-07 V_hig
+ 1.554010000e-07 V_hig
+ 1.555000000e-07 V_hig
+ 1.555010000e-07 V_hig
+ 1.556000000e-07 V_hig
+ 1.556010000e-07 V_hig
+ 1.557000000e-07 V_hig
+ 1.557010000e-07 V_hig
+ 1.558000000e-07 V_hig
+ 1.558010000e-07 V_hig
+ 1.559000000e-07 V_hig
+ 1.559010000e-07 V_hig
+ 1.560000000e-07 V_hig
+ 1.560010000e-07 V_hig
+ 1.561000000e-07 V_hig
+ 1.561010000e-07 V_hig
+ 1.562000000e-07 V_hig
+ 1.562010000e-07 V_hig
+ 1.563000000e-07 V_hig
+ 1.563010000e-07 V_hig
+ 1.564000000e-07 V_hig
+ 1.564010000e-07 V_hig
+ 1.565000000e-07 V_hig
+ 1.565010000e-07 V_hig
+ 1.566000000e-07 V_hig
+ 1.566010000e-07 V_hig
+ 1.567000000e-07 V_hig
+ 1.567010000e-07 V_hig
+ 1.568000000e-07 V_hig
+ 1.568010000e-07 V_hig
+ 1.569000000e-07 V_hig
+ 1.569010000e-07 V_low
+ 1.570000000e-07 V_low
+ 1.570010000e-07 V_low
+ 1.571000000e-07 V_low
+ 1.571010000e-07 V_low
+ 1.572000000e-07 V_low
+ 1.572010000e-07 V_low
+ 1.573000000e-07 V_low
+ 1.573010000e-07 V_low
+ 1.574000000e-07 V_low
+ 1.574010000e-07 V_low
+ 1.575000000e-07 V_low
+ 1.575010000e-07 V_low
+ 1.576000000e-07 V_low
+ 1.576010000e-07 V_low
+ 1.577000000e-07 V_low
+ 1.577010000e-07 V_low
+ 1.578000000e-07 V_low
+ 1.578010000e-07 V_low
+ 1.579000000e-07 V_low
+ 1.579010000e-07 V_hig
+ 1.580000000e-07 V_hig
+ 1.580010000e-07 V_hig
+ 1.581000000e-07 V_hig
+ 1.581010000e-07 V_hig
+ 1.582000000e-07 V_hig
+ 1.582010000e-07 V_hig
+ 1.583000000e-07 V_hig
+ 1.583010000e-07 V_hig
+ 1.584000000e-07 V_hig
+ 1.584010000e-07 V_hig
+ 1.585000000e-07 V_hig
+ 1.585010000e-07 V_hig
+ 1.586000000e-07 V_hig
+ 1.586010000e-07 V_hig
+ 1.587000000e-07 V_hig
+ 1.587010000e-07 V_hig
+ 1.588000000e-07 V_hig
+ 1.588010000e-07 V_hig
+ 1.589000000e-07 V_hig
+ 1.589010000e-07 V_hig
+ 1.590000000e-07 V_hig
+ 1.590010000e-07 V_hig
+ 1.591000000e-07 V_hig
+ 1.591010000e-07 V_hig
+ 1.592000000e-07 V_hig
+ 1.592010000e-07 V_hig
+ 1.593000000e-07 V_hig
+ 1.593010000e-07 V_hig
+ 1.594000000e-07 V_hig
+ 1.594010000e-07 V_hig
+ 1.595000000e-07 V_hig
+ 1.595010000e-07 V_hig
+ 1.596000000e-07 V_hig
+ 1.596010000e-07 V_hig
+ 1.597000000e-07 V_hig
+ 1.597010000e-07 V_hig
+ 1.598000000e-07 V_hig
+ 1.598010000e-07 V_hig
+ 1.599000000e-07 V_hig
+ 1.599010000e-07 V_low
+ 1.600000000e-07 V_low
+ 1.600010000e-07 V_low
+ 1.601000000e-07 V_low
+ 1.601010000e-07 V_low
+ 1.602000000e-07 V_low
+ 1.602010000e-07 V_low
+ 1.603000000e-07 V_low
+ 1.603010000e-07 V_low
+ 1.604000000e-07 V_low
+ 1.604010000e-07 V_low
+ 1.605000000e-07 V_low
+ 1.605010000e-07 V_low
+ 1.606000000e-07 V_low
+ 1.606010000e-07 V_low
+ 1.607000000e-07 V_low
+ 1.607010000e-07 V_low
+ 1.608000000e-07 V_low
+ 1.608010000e-07 V_low
+ 1.609000000e-07 V_low
+ 1.609010000e-07 V_low
+ 1.610000000e-07 V_low
+ 1.610010000e-07 V_low
+ 1.611000000e-07 V_low
+ 1.611010000e-07 V_low
+ 1.612000000e-07 V_low
+ 1.612010000e-07 V_low
+ 1.613000000e-07 V_low
+ 1.613010000e-07 V_low
+ 1.614000000e-07 V_low
+ 1.614010000e-07 V_low
+ 1.615000000e-07 V_low
+ 1.615010000e-07 V_low
+ 1.616000000e-07 V_low
+ 1.616010000e-07 V_low
+ 1.617000000e-07 V_low
+ 1.617010000e-07 V_low
+ 1.618000000e-07 V_low
+ 1.618010000e-07 V_low
+ 1.619000000e-07 V_low
+ 1.619010000e-07 V_low
+ 1.620000000e-07 V_low
+ 1.620010000e-07 V_low
+ 1.621000000e-07 V_low
+ 1.621010000e-07 V_low
+ 1.622000000e-07 V_low
+ 1.622010000e-07 V_low
+ 1.623000000e-07 V_low
+ 1.623010000e-07 V_low
+ 1.624000000e-07 V_low
+ 1.624010000e-07 V_low
+ 1.625000000e-07 V_low
+ 1.625010000e-07 V_low
+ 1.626000000e-07 V_low
+ 1.626010000e-07 V_low
+ 1.627000000e-07 V_low
+ 1.627010000e-07 V_low
+ 1.628000000e-07 V_low
+ 1.628010000e-07 V_low
+ 1.629000000e-07 V_low
+ 1.629010000e-07 V_low
+ 1.630000000e-07 V_low
+ 1.630010000e-07 V_low
+ 1.631000000e-07 V_low
+ 1.631010000e-07 V_low
+ 1.632000000e-07 V_low
+ 1.632010000e-07 V_low
+ 1.633000000e-07 V_low
+ 1.633010000e-07 V_low
+ 1.634000000e-07 V_low
+ 1.634010000e-07 V_low
+ 1.635000000e-07 V_low
+ 1.635010000e-07 V_low
+ 1.636000000e-07 V_low
+ 1.636010000e-07 V_low
+ 1.637000000e-07 V_low
+ 1.637010000e-07 V_low
+ 1.638000000e-07 V_low
+ 1.638010000e-07 V_low
+ 1.639000000e-07 V_low
+ 1.639010000e-07 V_low
+ 1.640000000e-07 V_low
+ 1.640010000e-07 V_low
+ 1.641000000e-07 V_low
+ 1.641010000e-07 V_low
+ 1.642000000e-07 V_low
+ 1.642010000e-07 V_low
+ 1.643000000e-07 V_low
+ 1.643010000e-07 V_low
+ 1.644000000e-07 V_low
+ 1.644010000e-07 V_low
+ 1.645000000e-07 V_low
+ 1.645010000e-07 V_low
+ 1.646000000e-07 V_low
+ 1.646010000e-07 V_low
+ 1.647000000e-07 V_low
+ 1.647010000e-07 V_low
+ 1.648000000e-07 V_low
+ 1.648010000e-07 V_low
+ 1.649000000e-07 V_low
+ 1.649010000e-07 V_hig
+ 1.650000000e-07 V_hig
+ 1.650010000e-07 V_hig
+ 1.651000000e-07 V_hig
+ 1.651010000e-07 V_hig
+ 1.652000000e-07 V_hig
+ 1.652010000e-07 V_hig
+ 1.653000000e-07 V_hig
+ 1.653010000e-07 V_hig
+ 1.654000000e-07 V_hig
+ 1.654010000e-07 V_hig
+ 1.655000000e-07 V_hig
+ 1.655010000e-07 V_hig
+ 1.656000000e-07 V_hig
+ 1.656010000e-07 V_hig
+ 1.657000000e-07 V_hig
+ 1.657010000e-07 V_hig
+ 1.658000000e-07 V_hig
+ 1.658010000e-07 V_hig
+ 1.659000000e-07 V_hig
+ 1.659010000e-07 V_low
+ 1.660000000e-07 V_low
+ 1.660010000e-07 V_low
+ 1.661000000e-07 V_low
+ 1.661010000e-07 V_low
+ 1.662000000e-07 V_low
+ 1.662010000e-07 V_low
+ 1.663000000e-07 V_low
+ 1.663010000e-07 V_low
+ 1.664000000e-07 V_low
+ 1.664010000e-07 V_low
+ 1.665000000e-07 V_low
+ 1.665010000e-07 V_low
+ 1.666000000e-07 V_low
+ 1.666010000e-07 V_low
+ 1.667000000e-07 V_low
+ 1.667010000e-07 V_low
+ 1.668000000e-07 V_low
+ 1.668010000e-07 V_low
+ 1.669000000e-07 V_low
+ 1.669010000e-07 V_hig
+ 1.670000000e-07 V_hig
+ 1.670010000e-07 V_hig
+ 1.671000000e-07 V_hig
+ 1.671010000e-07 V_hig
+ 1.672000000e-07 V_hig
+ 1.672010000e-07 V_hig
+ 1.673000000e-07 V_hig
+ 1.673010000e-07 V_hig
+ 1.674000000e-07 V_hig
+ 1.674010000e-07 V_hig
+ 1.675000000e-07 V_hig
+ 1.675010000e-07 V_hig
+ 1.676000000e-07 V_hig
+ 1.676010000e-07 V_hig
+ 1.677000000e-07 V_hig
+ 1.677010000e-07 V_hig
+ 1.678000000e-07 V_hig
+ 1.678010000e-07 V_hig
+ 1.679000000e-07 V_hig
+ 1.679010000e-07 V_hig
+ 1.680000000e-07 V_hig
+ 1.680010000e-07 V_hig
+ 1.681000000e-07 V_hig
+ 1.681010000e-07 V_hig
+ 1.682000000e-07 V_hig
+ 1.682010000e-07 V_hig
+ 1.683000000e-07 V_hig
+ 1.683010000e-07 V_hig
+ 1.684000000e-07 V_hig
+ 1.684010000e-07 V_hig
+ 1.685000000e-07 V_hig
+ 1.685010000e-07 V_hig
+ 1.686000000e-07 V_hig
+ 1.686010000e-07 V_hig
+ 1.687000000e-07 V_hig
+ 1.687010000e-07 V_hig
+ 1.688000000e-07 V_hig
+ 1.688010000e-07 V_hig
+ 1.689000000e-07 V_hig
+ 1.689010000e-07 V_hig
+ 1.690000000e-07 V_hig
+ 1.690010000e-07 V_hig
+ 1.691000000e-07 V_hig
+ 1.691010000e-07 V_hig
+ 1.692000000e-07 V_hig
+ 1.692010000e-07 V_hig
+ 1.693000000e-07 V_hig
+ 1.693010000e-07 V_hig
+ 1.694000000e-07 V_hig
+ 1.694010000e-07 V_hig
+ 1.695000000e-07 V_hig
+ 1.695010000e-07 V_hig
+ 1.696000000e-07 V_hig
+ 1.696010000e-07 V_hig
+ 1.697000000e-07 V_hig
+ 1.697010000e-07 V_hig
+ 1.698000000e-07 V_hig
+ 1.698010000e-07 V_hig
+ 1.699000000e-07 V_hig
+ 1.699010000e-07 V_hig
+ 1.700000000e-07 V_hig
+ 1.700010000e-07 V_hig
+ 1.701000000e-07 V_hig
+ 1.701010000e-07 V_hig
+ 1.702000000e-07 V_hig
+ 1.702010000e-07 V_hig
+ 1.703000000e-07 V_hig
+ 1.703010000e-07 V_hig
+ 1.704000000e-07 V_hig
+ 1.704010000e-07 V_hig
+ 1.705000000e-07 V_hig
+ 1.705010000e-07 V_hig
+ 1.706000000e-07 V_hig
+ 1.706010000e-07 V_hig
+ 1.707000000e-07 V_hig
+ 1.707010000e-07 V_hig
+ 1.708000000e-07 V_hig
+ 1.708010000e-07 V_hig
+ 1.709000000e-07 V_hig
+ 1.709010000e-07 V_hig
+ 1.710000000e-07 V_hig
+ 1.710010000e-07 V_hig
+ 1.711000000e-07 V_hig
+ 1.711010000e-07 V_hig
+ 1.712000000e-07 V_hig
+ 1.712010000e-07 V_hig
+ 1.713000000e-07 V_hig
+ 1.713010000e-07 V_hig
+ 1.714000000e-07 V_hig
+ 1.714010000e-07 V_hig
+ 1.715000000e-07 V_hig
+ 1.715010000e-07 V_hig
+ 1.716000000e-07 V_hig
+ 1.716010000e-07 V_hig
+ 1.717000000e-07 V_hig
+ 1.717010000e-07 V_hig
+ 1.718000000e-07 V_hig
+ 1.718010000e-07 V_hig
+ 1.719000000e-07 V_hig
+ 1.719010000e-07 V_low
+ 1.720000000e-07 V_low
+ 1.720010000e-07 V_low
+ 1.721000000e-07 V_low
+ 1.721010000e-07 V_low
+ 1.722000000e-07 V_low
+ 1.722010000e-07 V_low
+ 1.723000000e-07 V_low
+ 1.723010000e-07 V_low
+ 1.724000000e-07 V_low
+ 1.724010000e-07 V_low
+ 1.725000000e-07 V_low
+ 1.725010000e-07 V_low
+ 1.726000000e-07 V_low
+ 1.726010000e-07 V_low
+ 1.727000000e-07 V_low
+ 1.727010000e-07 V_low
+ 1.728000000e-07 V_low
+ 1.728010000e-07 V_low
+ 1.729000000e-07 V_low
+ 1.729010000e-07 V_hig
+ 1.730000000e-07 V_hig
+ 1.730010000e-07 V_hig
+ 1.731000000e-07 V_hig
+ 1.731010000e-07 V_hig
+ 1.732000000e-07 V_hig
+ 1.732010000e-07 V_hig
+ 1.733000000e-07 V_hig
+ 1.733010000e-07 V_hig
+ 1.734000000e-07 V_hig
+ 1.734010000e-07 V_hig
+ 1.735000000e-07 V_hig
+ 1.735010000e-07 V_hig
+ 1.736000000e-07 V_hig
+ 1.736010000e-07 V_hig
+ 1.737000000e-07 V_hig
+ 1.737010000e-07 V_hig
+ 1.738000000e-07 V_hig
+ 1.738010000e-07 V_hig
+ 1.739000000e-07 V_hig
+ 1.739010000e-07 V_hig
+ 1.740000000e-07 V_hig
+ 1.740010000e-07 V_hig
+ 1.741000000e-07 V_hig
+ 1.741010000e-07 V_hig
+ 1.742000000e-07 V_hig
+ 1.742010000e-07 V_hig
+ 1.743000000e-07 V_hig
+ 1.743010000e-07 V_hig
+ 1.744000000e-07 V_hig
+ 1.744010000e-07 V_hig
+ 1.745000000e-07 V_hig
+ 1.745010000e-07 V_hig
+ 1.746000000e-07 V_hig
+ 1.746010000e-07 V_hig
+ 1.747000000e-07 V_hig
+ 1.747010000e-07 V_hig
+ 1.748000000e-07 V_hig
+ 1.748010000e-07 V_hig
+ 1.749000000e-07 V_hig
+ 1.749010000e-07 V_hig
+ 1.750000000e-07 V_hig
+ 1.750010000e-07 V_hig
+ 1.751000000e-07 V_hig
+ 1.751010000e-07 V_hig
+ 1.752000000e-07 V_hig
+ 1.752010000e-07 V_hig
+ 1.753000000e-07 V_hig
+ 1.753010000e-07 V_hig
+ 1.754000000e-07 V_hig
+ 1.754010000e-07 V_hig
+ 1.755000000e-07 V_hig
+ 1.755010000e-07 V_hig
+ 1.756000000e-07 V_hig
+ 1.756010000e-07 V_hig
+ 1.757000000e-07 V_hig
+ 1.757010000e-07 V_hig
+ 1.758000000e-07 V_hig
+ 1.758010000e-07 V_hig
+ 1.759000000e-07 V_hig
+ 1.759010000e-07 V_low
+ 1.760000000e-07 V_low
+ 1.760010000e-07 V_low
+ 1.761000000e-07 V_low
+ 1.761010000e-07 V_low
+ 1.762000000e-07 V_low
+ 1.762010000e-07 V_low
+ 1.763000000e-07 V_low
+ 1.763010000e-07 V_low
+ 1.764000000e-07 V_low
+ 1.764010000e-07 V_low
+ 1.765000000e-07 V_low
+ 1.765010000e-07 V_low
+ 1.766000000e-07 V_low
+ 1.766010000e-07 V_low
+ 1.767000000e-07 V_low
+ 1.767010000e-07 V_low
+ 1.768000000e-07 V_low
+ 1.768010000e-07 V_low
+ 1.769000000e-07 V_low
+ 1.769010000e-07 V_hig
+ 1.770000000e-07 V_hig
+ 1.770010000e-07 V_hig
+ 1.771000000e-07 V_hig
+ 1.771010000e-07 V_hig
+ 1.772000000e-07 V_hig
+ 1.772010000e-07 V_hig
+ 1.773000000e-07 V_hig
+ 1.773010000e-07 V_hig
+ 1.774000000e-07 V_hig
+ 1.774010000e-07 V_hig
+ 1.775000000e-07 V_hig
+ 1.775010000e-07 V_hig
+ 1.776000000e-07 V_hig
+ 1.776010000e-07 V_hig
+ 1.777000000e-07 V_hig
+ 1.777010000e-07 V_hig
+ 1.778000000e-07 V_hig
+ 1.778010000e-07 V_hig
+ 1.779000000e-07 V_hig
+ 1.779010000e-07 V_hig
+ 1.780000000e-07 V_hig
+ 1.780010000e-07 V_hig
+ 1.781000000e-07 V_hig
+ 1.781010000e-07 V_hig
+ 1.782000000e-07 V_hig
+ 1.782010000e-07 V_hig
+ 1.783000000e-07 V_hig
+ 1.783010000e-07 V_hig
+ 1.784000000e-07 V_hig
+ 1.784010000e-07 V_hig
+ 1.785000000e-07 V_hig
+ 1.785010000e-07 V_hig
+ 1.786000000e-07 V_hig
+ 1.786010000e-07 V_hig
+ 1.787000000e-07 V_hig
+ 1.787010000e-07 V_hig
+ 1.788000000e-07 V_hig
+ 1.788010000e-07 V_hig
+ 1.789000000e-07 V_hig
+ 1.789010000e-07 V_low
+ 1.790000000e-07 V_low
+ 1.790010000e-07 V_low
+ 1.791000000e-07 V_low
+ 1.791010000e-07 V_low
+ 1.792000000e-07 V_low
+ 1.792010000e-07 V_low
+ 1.793000000e-07 V_low
+ 1.793010000e-07 V_low
+ 1.794000000e-07 V_low
+ 1.794010000e-07 V_low
+ 1.795000000e-07 V_low
+ 1.795010000e-07 V_low
+ 1.796000000e-07 V_low
+ 1.796010000e-07 V_low
+ 1.797000000e-07 V_low
+ 1.797010000e-07 V_low
+ 1.798000000e-07 V_low
+ 1.798010000e-07 V_low
+ 1.799000000e-07 V_low
+ 1.799010000e-07 V_hig
+ 1.800000000e-07 V_hig
+ 1.800010000e-07 V_hig
+ 1.801000000e-07 V_hig
+ 1.801010000e-07 V_hig
+ 1.802000000e-07 V_hig
+ 1.802010000e-07 V_hig
+ 1.803000000e-07 V_hig
+ 1.803010000e-07 V_hig
+ 1.804000000e-07 V_hig
+ 1.804010000e-07 V_hig
+ 1.805000000e-07 V_hig
+ 1.805010000e-07 V_hig
+ 1.806000000e-07 V_hig
+ 1.806010000e-07 V_hig
+ 1.807000000e-07 V_hig
+ 1.807010000e-07 V_hig
+ 1.808000000e-07 V_hig
+ 1.808010000e-07 V_hig
+ 1.809000000e-07 V_hig
+ 1.809010000e-07 V_hig
+ 1.810000000e-07 V_hig
+ 1.810010000e-07 V_hig
+ 1.811000000e-07 V_hig
+ 1.811010000e-07 V_hig
+ 1.812000000e-07 V_hig
+ 1.812010000e-07 V_hig
+ 1.813000000e-07 V_hig
+ 1.813010000e-07 V_hig
+ 1.814000000e-07 V_hig
+ 1.814010000e-07 V_hig
+ 1.815000000e-07 V_hig
+ 1.815010000e-07 V_hig
+ 1.816000000e-07 V_hig
+ 1.816010000e-07 V_hig
+ 1.817000000e-07 V_hig
+ 1.817010000e-07 V_hig
+ 1.818000000e-07 V_hig
+ 1.818010000e-07 V_hig
+ 1.819000000e-07 V_hig
+ 1.819010000e-07 V_low
+ 1.820000000e-07 V_low
+ 1.820010000e-07 V_low
+ 1.821000000e-07 V_low
+ 1.821010000e-07 V_low
+ 1.822000000e-07 V_low
+ 1.822010000e-07 V_low
+ 1.823000000e-07 V_low
+ 1.823010000e-07 V_low
+ 1.824000000e-07 V_low
+ 1.824010000e-07 V_low
+ 1.825000000e-07 V_low
+ 1.825010000e-07 V_low
+ 1.826000000e-07 V_low
+ 1.826010000e-07 V_low
+ 1.827000000e-07 V_low
+ 1.827010000e-07 V_low
+ 1.828000000e-07 V_low
+ 1.828010000e-07 V_low
+ 1.829000000e-07 V_low
+ 1.829010000e-07 V_hig
+ 1.830000000e-07 V_hig
+ 1.830010000e-07 V_hig
+ 1.831000000e-07 V_hig
+ 1.831010000e-07 V_hig
+ 1.832000000e-07 V_hig
+ 1.832010000e-07 V_hig
+ 1.833000000e-07 V_hig
+ 1.833010000e-07 V_hig
+ 1.834000000e-07 V_hig
+ 1.834010000e-07 V_hig
+ 1.835000000e-07 V_hig
+ 1.835010000e-07 V_hig
+ 1.836000000e-07 V_hig
+ 1.836010000e-07 V_hig
+ 1.837000000e-07 V_hig
+ 1.837010000e-07 V_hig
+ 1.838000000e-07 V_hig
+ 1.838010000e-07 V_hig
+ 1.839000000e-07 V_hig
+ 1.839010000e-07 V_low
+ 1.840000000e-07 V_low
+ 1.840010000e-07 V_low
+ 1.841000000e-07 V_low
+ 1.841010000e-07 V_low
+ 1.842000000e-07 V_low
+ 1.842010000e-07 V_low
+ 1.843000000e-07 V_low
+ 1.843010000e-07 V_low
+ 1.844000000e-07 V_low
+ 1.844010000e-07 V_low
+ 1.845000000e-07 V_low
+ 1.845010000e-07 V_low
+ 1.846000000e-07 V_low
+ 1.846010000e-07 V_low
+ 1.847000000e-07 V_low
+ 1.847010000e-07 V_low
+ 1.848000000e-07 V_low
+ 1.848010000e-07 V_low
+ 1.849000000e-07 V_low
+ 1.849010000e-07 V_hig
+ 1.850000000e-07 V_hig
+ 1.850010000e-07 V_hig
+ 1.851000000e-07 V_hig
+ 1.851010000e-07 V_hig
+ 1.852000000e-07 V_hig
+ 1.852010000e-07 V_hig
+ 1.853000000e-07 V_hig
+ 1.853010000e-07 V_hig
+ 1.854000000e-07 V_hig
+ 1.854010000e-07 V_hig
+ 1.855000000e-07 V_hig
+ 1.855010000e-07 V_hig
+ 1.856000000e-07 V_hig
+ 1.856010000e-07 V_hig
+ 1.857000000e-07 V_hig
+ 1.857010000e-07 V_hig
+ 1.858000000e-07 V_hig
+ 1.858010000e-07 V_hig
+ 1.859000000e-07 V_hig
+ 1.859010000e-07 V_hig
+ 1.860000000e-07 V_hig
+ 1.860010000e-07 V_hig
+ 1.861000000e-07 V_hig
+ 1.861010000e-07 V_hig
+ 1.862000000e-07 V_hig
+ 1.862010000e-07 V_hig
+ 1.863000000e-07 V_hig
+ 1.863010000e-07 V_hig
+ 1.864000000e-07 V_hig
+ 1.864010000e-07 V_hig
+ 1.865000000e-07 V_hig
+ 1.865010000e-07 V_hig
+ 1.866000000e-07 V_hig
+ 1.866010000e-07 V_hig
+ 1.867000000e-07 V_hig
+ 1.867010000e-07 V_hig
+ 1.868000000e-07 V_hig
+ 1.868010000e-07 V_hig
+ 1.869000000e-07 V_hig
+ 1.869010000e-07 V_hig
+ 1.870000000e-07 V_hig
+ 1.870010000e-07 V_hig
+ 1.871000000e-07 V_hig
+ 1.871010000e-07 V_hig
+ 1.872000000e-07 V_hig
+ 1.872010000e-07 V_hig
+ 1.873000000e-07 V_hig
+ 1.873010000e-07 V_hig
+ 1.874000000e-07 V_hig
+ 1.874010000e-07 V_hig
+ 1.875000000e-07 V_hig
+ 1.875010000e-07 V_hig
+ 1.876000000e-07 V_hig
+ 1.876010000e-07 V_hig
+ 1.877000000e-07 V_hig
+ 1.877010000e-07 V_hig
+ 1.878000000e-07 V_hig
+ 1.878010000e-07 V_hig
+ 1.879000000e-07 V_hig
+ 1.879010000e-07 V_low
+ 1.880000000e-07 V_low
+ 1.880010000e-07 V_low
+ 1.881000000e-07 V_low
+ 1.881010000e-07 V_low
+ 1.882000000e-07 V_low
+ 1.882010000e-07 V_low
+ 1.883000000e-07 V_low
+ 1.883010000e-07 V_low
+ 1.884000000e-07 V_low
+ 1.884010000e-07 V_low
+ 1.885000000e-07 V_low
+ 1.885010000e-07 V_low
+ 1.886000000e-07 V_low
+ 1.886010000e-07 V_low
+ 1.887000000e-07 V_low
+ 1.887010000e-07 V_low
+ 1.888000000e-07 V_low
+ 1.888010000e-07 V_low
+ 1.889000000e-07 V_low
+ 1.889010000e-07 V_low
+ 1.890000000e-07 V_low
+ 1.890010000e-07 V_low
+ 1.891000000e-07 V_low
+ 1.891010000e-07 V_low
+ 1.892000000e-07 V_low
+ 1.892010000e-07 V_low
+ 1.893000000e-07 V_low
+ 1.893010000e-07 V_low
+ 1.894000000e-07 V_low
+ 1.894010000e-07 V_low
+ 1.895000000e-07 V_low
+ 1.895010000e-07 V_low
+ 1.896000000e-07 V_low
+ 1.896010000e-07 V_low
+ 1.897000000e-07 V_low
+ 1.897010000e-07 V_low
+ 1.898000000e-07 V_low
+ 1.898010000e-07 V_low
+ 1.899000000e-07 V_low
+ 1.899010000e-07 V_hig
+ 1.900000000e-07 V_hig
+ 1.900010000e-07 V_hig
+ 1.901000000e-07 V_hig
+ 1.901010000e-07 V_hig
+ 1.902000000e-07 V_hig
+ 1.902010000e-07 V_hig
+ 1.903000000e-07 V_hig
+ 1.903010000e-07 V_hig
+ 1.904000000e-07 V_hig
+ 1.904010000e-07 V_hig
+ 1.905000000e-07 V_hig
+ 1.905010000e-07 V_hig
+ 1.906000000e-07 V_hig
+ 1.906010000e-07 V_hig
+ 1.907000000e-07 V_hig
+ 1.907010000e-07 V_hig
+ 1.908000000e-07 V_hig
+ 1.908010000e-07 V_hig
+ 1.909000000e-07 V_hig
+ 1.909010000e-07 V_low
+ 1.910000000e-07 V_low
+ 1.910010000e-07 V_low
+ 1.911000000e-07 V_low
+ 1.911010000e-07 V_low
+ 1.912000000e-07 V_low
+ 1.912010000e-07 V_low
+ 1.913000000e-07 V_low
+ 1.913010000e-07 V_low
+ 1.914000000e-07 V_low
+ 1.914010000e-07 V_low
+ 1.915000000e-07 V_low
+ 1.915010000e-07 V_low
+ 1.916000000e-07 V_low
+ 1.916010000e-07 V_low
+ 1.917000000e-07 V_low
+ 1.917010000e-07 V_low
+ 1.918000000e-07 V_low
+ 1.918010000e-07 V_low
+ 1.919000000e-07 V_low
+ 1.919010000e-07 V_low
+ 1.920000000e-07 V_low
+ 1.920010000e-07 V_low
+ 1.921000000e-07 V_low
+ 1.921010000e-07 V_low
+ 1.922000000e-07 V_low
+ 1.922010000e-07 V_low
+ 1.923000000e-07 V_low
+ 1.923010000e-07 V_low
+ 1.924000000e-07 V_low
+ 1.924010000e-07 V_low
+ 1.925000000e-07 V_low
+ 1.925010000e-07 V_low
+ 1.926000000e-07 V_low
+ 1.926010000e-07 V_low
+ 1.927000000e-07 V_low
+ 1.927010000e-07 V_low
+ 1.928000000e-07 V_low
+ 1.928010000e-07 V_low
+ 1.929000000e-07 V_low
+ 1.929010000e-07 V_hig
+ 1.930000000e-07 V_hig
+ 1.930010000e-07 V_hig
+ 1.931000000e-07 V_hig
+ 1.931010000e-07 V_hig
+ 1.932000000e-07 V_hig
+ 1.932010000e-07 V_hig
+ 1.933000000e-07 V_hig
+ 1.933010000e-07 V_hig
+ 1.934000000e-07 V_hig
+ 1.934010000e-07 V_hig
+ 1.935000000e-07 V_hig
+ 1.935010000e-07 V_hig
+ 1.936000000e-07 V_hig
+ 1.936010000e-07 V_hig
+ 1.937000000e-07 V_hig
+ 1.937010000e-07 V_hig
+ 1.938000000e-07 V_hig
+ 1.938010000e-07 V_hig
+ 1.939000000e-07 V_hig
+ 1.939010000e-07 V_hig
+ 1.940000000e-07 V_hig
+ 1.940010000e-07 V_hig
+ 1.941000000e-07 V_hig
+ 1.941010000e-07 V_hig
+ 1.942000000e-07 V_hig
+ 1.942010000e-07 V_hig
+ 1.943000000e-07 V_hig
+ 1.943010000e-07 V_hig
+ 1.944000000e-07 V_hig
+ 1.944010000e-07 V_hig
+ 1.945000000e-07 V_hig
+ 1.945010000e-07 V_hig
+ 1.946000000e-07 V_hig
+ 1.946010000e-07 V_hig
+ 1.947000000e-07 V_hig
+ 1.947010000e-07 V_hig
+ 1.948000000e-07 V_hig
+ 1.948010000e-07 V_hig
+ 1.949000000e-07 V_hig
+ 1.949010000e-07 V_low
+ 1.950000000e-07 V_low
+ 1.950010000e-07 V_low
+ 1.951000000e-07 V_low
+ 1.951010000e-07 V_low
+ 1.952000000e-07 V_low
+ 1.952010000e-07 V_low
+ 1.953000000e-07 V_low
+ 1.953010000e-07 V_low
+ 1.954000000e-07 V_low
+ 1.954010000e-07 V_low
+ 1.955000000e-07 V_low
+ 1.955010000e-07 V_low
+ 1.956000000e-07 V_low
+ 1.956010000e-07 V_low
+ 1.957000000e-07 V_low
+ 1.957010000e-07 V_low
+ 1.958000000e-07 V_low
+ 1.958010000e-07 V_low
+ 1.959000000e-07 V_low
+ 1.959010000e-07 V_low
+ 1.960000000e-07 V_low
+ 1.960010000e-07 V_low
+ 1.961000000e-07 V_low
+ 1.961010000e-07 V_low
+ 1.962000000e-07 V_low
+ 1.962010000e-07 V_low
+ 1.963000000e-07 V_low
+ 1.963010000e-07 V_low
+ 1.964000000e-07 V_low
+ 1.964010000e-07 V_low
+ 1.965000000e-07 V_low
+ 1.965010000e-07 V_low
+ 1.966000000e-07 V_low
+ 1.966010000e-07 V_low
+ 1.967000000e-07 V_low
+ 1.967010000e-07 V_low
+ 1.968000000e-07 V_low
+ 1.968010000e-07 V_low
+ 1.969000000e-07 V_low
+ 1.969010000e-07 V_hig
+ 1.970000000e-07 V_hig
+ 1.970010000e-07 V_hig
+ 1.971000000e-07 V_hig
+ 1.971010000e-07 V_hig
+ 1.972000000e-07 V_hig
+ 1.972010000e-07 V_hig
+ 1.973000000e-07 V_hig
+ 1.973010000e-07 V_hig
+ 1.974000000e-07 V_hig
+ 1.974010000e-07 V_hig
+ 1.975000000e-07 V_hig
+ 1.975010000e-07 V_hig
+ 1.976000000e-07 V_hig
+ 1.976010000e-07 V_hig
+ 1.977000000e-07 V_hig
+ 1.977010000e-07 V_hig
+ 1.978000000e-07 V_hig
+ 1.978010000e-07 V_hig
+ 1.979000000e-07 V_hig
+ 1.979010000e-07 V_hig
+ 1.980000000e-07 V_hig
+ 1.980010000e-07 V_hig
+ 1.981000000e-07 V_hig
+ 1.981010000e-07 V_hig
+ 1.982000000e-07 V_hig
+ 1.982010000e-07 V_hig
+ 1.983000000e-07 V_hig
+ 1.983010000e-07 V_hig
+ 1.984000000e-07 V_hig
+ 1.984010000e-07 V_hig
+ 1.985000000e-07 V_hig
+ 1.985010000e-07 V_hig
+ 1.986000000e-07 V_hig
+ 1.986010000e-07 V_hig
+ 1.987000000e-07 V_hig
+ 1.987010000e-07 V_hig
+ 1.988000000e-07 V_hig
+ 1.988010000e-07 V_hig
+ 1.989000000e-07 V_hig
+ 1.989010000e-07 V_low
+ 1.990000000e-07 V_low
+ 1.990010000e-07 V_low
+ 1.991000000e-07 V_low
+ 1.991010000e-07 V_low
+ 1.992000000e-07 V_low
+ 1.992010000e-07 V_low
+ 1.993000000e-07 V_low
+ 1.993010000e-07 V_low
+ 1.994000000e-07 V_low
+ 1.994010000e-07 V_low
+ 1.995000000e-07 V_low
+ 1.995010000e-07 V_low
+ 1.996000000e-07 V_low
+ 1.996010000e-07 V_low
+ 1.997000000e-07 V_low
+ 1.997010000e-07 V_low
+ 1.998000000e-07 V_low
+ 1.998010000e-07 V_low
+ 1.999000000e-07 V_low
+ 1.999010000e-07 V_hig
+ 2.000000000e-07 V_hig
+ 2.000010000e-07 V_hig
+ 2.001000000e-07 V_hig
+ 2.001010000e-07 V_hig
+ 2.002000000e-07 V_hig
+ 2.002010000e-07 V_hig
+ 2.003000000e-07 V_hig
+ 2.003010000e-07 V_hig
+ 2.004000000e-07 V_hig
+ 2.004010000e-07 V_hig
+ 2.005000000e-07 V_hig
+ 2.005010000e-07 V_hig
+ 2.006000000e-07 V_hig
+ 2.006010000e-07 V_hig
+ 2.007000000e-07 V_hig
+ 2.007010000e-07 V_hig
+ 2.008000000e-07 V_hig
+ 2.008010000e-07 V_hig
+ 2.009000000e-07 V_hig
+ 2.009010000e-07 V_hig
+ 2.010000000e-07 V_hig
+ 2.010010000e-07 V_hig
+ 2.011000000e-07 V_hig
+ 2.011010000e-07 V_hig
+ 2.012000000e-07 V_hig
+ 2.012010000e-07 V_hig
+ 2.013000000e-07 V_hig
+ 2.013010000e-07 V_hig
+ 2.014000000e-07 V_hig
+ 2.014010000e-07 V_hig
+ 2.015000000e-07 V_hig
+ 2.015010000e-07 V_hig
+ 2.016000000e-07 V_hig
+ 2.016010000e-07 V_hig
+ 2.017000000e-07 V_hig
+ 2.017010000e-07 V_hig
+ 2.018000000e-07 V_hig
+ 2.018010000e-07 V_hig
+ 2.019000000e-07 V_hig
+ 2.019010000e-07 V_low
+ 2.020000000e-07 V_low
+ 2.020010000e-07 V_low
+ 2.021000000e-07 V_low
+ 2.021010000e-07 V_low
+ 2.022000000e-07 V_low
+ 2.022010000e-07 V_low
+ 2.023000000e-07 V_low
+ 2.023010000e-07 V_low
+ 2.024000000e-07 V_low
+ 2.024010000e-07 V_low
+ 2.025000000e-07 V_low
+ 2.025010000e-07 V_low
+ 2.026000000e-07 V_low
+ 2.026010000e-07 V_low
+ 2.027000000e-07 V_low
+ 2.027010000e-07 V_low
+ 2.028000000e-07 V_low
+ 2.028010000e-07 V_low
+ 2.029000000e-07 V_low
+ 2.029010000e-07 V_low
+ 2.030000000e-07 V_low
+ 2.030010000e-07 V_low
+ 2.031000000e-07 V_low
+ 2.031010000e-07 V_low
+ 2.032000000e-07 V_low
+ 2.032010000e-07 V_low
+ 2.033000000e-07 V_low
+ 2.033010000e-07 V_low
+ 2.034000000e-07 V_low
+ 2.034010000e-07 V_low
+ 2.035000000e-07 V_low
+ 2.035010000e-07 V_low
+ 2.036000000e-07 V_low
+ 2.036010000e-07 V_low
+ 2.037000000e-07 V_low
+ 2.037010000e-07 V_low
+ 2.038000000e-07 V_low
+ 2.038010000e-07 V_low
+ 2.039000000e-07 V_low
+ 2.039010000e-07 V_low
+ 2.040000000e-07 V_low
+ 2.040010000e-07 V_low
+ 2.041000000e-07 V_low
+ 2.041010000e-07 V_low
+ 2.042000000e-07 V_low
+ 2.042010000e-07 V_low
+ 2.043000000e-07 V_low
+ 2.043010000e-07 V_low
+ 2.044000000e-07 V_low
+ 2.044010000e-07 V_low
+ 2.045000000e-07 V_low
+ 2.045010000e-07 V_low
+ 2.046000000e-07 V_low
+ 2.046010000e-07 V_low
+ 2.047000000e-07 V_low
+ 2.047010000e-07 V_low
+ 2.048000000e-07 V_low
+ 2.048010000e-07 V_low
+ 2.049000000e-07 V_low
+ 2.049010000e-07 V_low
+ 2.050000000e-07 V_low
+ 2.050010000e-07 V_low
+ 2.051000000e-07 V_low
+ 2.051010000e-07 V_low
+ 2.052000000e-07 V_low
+ 2.052010000e-07 V_low
+ 2.053000000e-07 V_low
+ 2.053010000e-07 V_low
+ 2.054000000e-07 V_low
+ 2.054010000e-07 V_low
+ 2.055000000e-07 V_low
+ 2.055010000e-07 V_low
+ 2.056000000e-07 V_low
+ 2.056010000e-07 V_low
+ 2.057000000e-07 V_low
+ 2.057010000e-07 V_low
+ 2.058000000e-07 V_low
+ 2.058010000e-07 V_low
+ 2.059000000e-07 V_low
+ 2.059010000e-07 V_low
+ 2.060000000e-07 V_low
+ 2.060010000e-07 V_low
+ 2.061000000e-07 V_low
+ 2.061010000e-07 V_low
+ 2.062000000e-07 V_low
+ 2.062010000e-07 V_low
+ 2.063000000e-07 V_low
+ 2.063010000e-07 V_low
+ 2.064000000e-07 V_low
+ 2.064010000e-07 V_low
+ 2.065000000e-07 V_low
+ 2.065010000e-07 V_low
+ 2.066000000e-07 V_low
+ 2.066010000e-07 V_low
+ 2.067000000e-07 V_low
+ 2.067010000e-07 V_low
+ 2.068000000e-07 V_low
+ 2.068010000e-07 V_low
+ 2.069000000e-07 V_low
+ 2.069010000e-07 V_low
+ 2.070000000e-07 V_low
+ 2.070010000e-07 V_low
+ 2.071000000e-07 V_low
+ 2.071010000e-07 V_low
+ 2.072000000e-07 V_low
+ 2.072010000e-07 V_low
+ 2.073000000e-07 V_low
+ 2.073010000e-07 V_low
+ 2.074000000e-07 V_low
+ 2.074010000e-07 V_low
+ 2.075000000e-07 V_low
+ 2.075010000e-07 V_low
+ 2.076000000e-07 V_low
+ 2.076010000e-07 V_low
+ 2.077000000e-07 V_low
+ 2.077010000e-07 V_low
+ 2.078000000e-07 V_low
+ 2.078010000e-07 V_low
+ 2.079000000e-07 V_low
+ 2.079010000e-07 V_hig
+ 2.080000000e-07 V_hig
+ 2.080010000e-07 V_hig
+ 2.081000000e-07 V_hig
+ 2.081010000e-07 V_hig
+ 2.082000000e-07 V_hig
+ 2.082010000e-07 V_hig
+ 2.083000000e-07 V_hig
+ 2.083010000e-07 V_hig
+ 2.084000000e-07 V_hig
+ 2.084010000e-07 V_hig
+ 2.085000000e-07 V_hig
+ 2.085010000e-07 V_hig
+ 2.086000000e-07 V_hig
+ 2.086010000e-07 V_hig
+ 2.087000000e-07 V_hig
+ 2.087010000e-07 V_hig
+ 2.088000000e-07 V_hig
+ 2.088010000e-07 V_hig
+ 2.089000000e-07 V_hig
+ 2.089010000e-07 V_low
+ 2.090000000e-07 V_low
+ 2.090010000e-07 V_low
+ 2.091000000e-07 V_low
+ 2.091010000e-07 V_low
+ 2.092000000e-07 V_low
+ 2.092010000e-07 V_low
+ 2.093000000e-07 V_low
+ 2.093010000e-07 V_low
+ 2.094000000e-07 V_low
+ 2.094010000e-07 V_low
+ 2.095000000e-07 V_low
+ 2.095010000e-07 V_low
+ 2.096000000e-07 V_low
+ 2.096010000e-07 V_low
+ 2.097000000e-07 V_low
+ 2.097010000e-07 V_low
+ 2.098000000e-07 V_low
+ 2.098010000e-07 V_low
+ 2.099000000e-07 V_low
+ 2.099010000e-07 V_low
+ 2.100000000e-07 V_low
+ 2.100010000e-07 V_low
+ 2.101000000e-07 V_low
+ 2.101010000e-07 V_low
+ 2.102000000e-07 V_low
+ 2.102010000e-07 V_low
+ 2.103000000e-07 V_low
+ 2.103010000e-07 V_low
+ 2.104000000e-07 V_low
+ 2.104010000e-07 V_low
+ 2.105000000e-07 V_low
+ 2.105010000e-07 V_low
+ 2.106000000e-07 V_low
+ 2.106010000e-07 V_low
+ 2.107000000e-07 V_low
+ 2.107010000e-07 V_low
+ 2.108000000e-07 V_low
+ 2.108010000e-07 V_low
+ 2.109000000e-07 V_low
+ 2.109010000e-07 V_hig
+ 2.110000000e-07 V_hig
+ 2.110010000e-07 V_hig
+ 2.111000000e-07 V_hig
+ 2.111010000e-07 V_hig
+ 2.112000000e-07 V_hig
+ 2.112010000e-07 V_hig
+ 2.113000000e-07 V_hig
+ 2.113010000e-07 V_hig
+ 2.114000000e-07 V_hig
+ 2.114010000e-07 V_hig
+ 2.115000000e-07 V_hig
+ 2.115010000e-07 V_hig
+ 2.116000000e-07 V_hig
+ 2.116010000e-07 V_hig
+ 2.117000000e-07 V_hig
+ 2.117010000e-07 V_hig
+ 2.118000000e-07 V_hig
+ 2.118010000e-07 V_hig
+ 2.119000000e-07 V_hig
+ 2.119010000e-07 V_low
+ 2.120000000e-07 V_low
+ 2.120010000e-07 V_low
+ 2.121000000e-07 V_low
+ 2.121010000e-07 V_low
+ 2.122000000e-07 V_low
+ 2.122010000e-07 V_low
+ 2.123000000e-07 V_low
+ 2.123010000e-07 V_low
+ 2.124000000e-07 V_low
+ 2.124010000e-07 V_low
+ 2.125000000e-07 V_low
+ 2.125010000e-07 V_low
+ 2.126000000e-07 V_low
+ 2.126010000e-07 V_low
+ 2.127000000e-07 V_low
+ 2.127010000e-07 V_low
+ 2.128000000e-07 V_low
+ 2.128010000e-07 V_low
+ 2.129000000e-07 V_low
+ 2.129010000e-07 V_low
+ 2.130000000e-07 V_low
+ 2.130010000e-07 V_low
+ 2.131000000e-07 V_low
+ 2.131010000e-07 V_low
+ 2.132000000e-07 V_low
+ 2.132010000e-07 V_low
+ 2.133000000e-07 V_low
+ 2.133010000e-07 V_low
+ 2.134000000e-07 V_low
+ 2.134010000e-07 V_low
+ 2.135000000e-07 V_low
+ 2.135010000e-07 V_low
+ 2.136000000e-07 V_low
+ 2.136010000e-07 V_low
+ 2.137000000e-07 V_low
+ 2.137010000e-07 V_low
+ 2.138000000e-07 V_low
+ 2.138010000e-07 V_low
+ 2.139000000e-07 V_low
+ 2.139010000e-07 V_low
+ 2.140000000e-07 V_low
+ 2.140010000e-07 V_low
+ 2.141000000e-07 V_low
+ 2.141010000e-07 V_low
+ 2.142000000e-07 V_low
+ 2.142010000e-07 V_low
+ 2.143000000e-07 V_low
+ 2.143010000e-07 V_low
+ 2.144000000e-07 V_low
+ 2.144010000e-07 V_low
+ 2.145000000e-07 V_low
+ 2.145010000e-07 V_low
+ 2.146000000e-07 V_low
+ 2.146010000e-07 V_low
+ 2.147000000e-07 V_low
+ 2.147010000e-07 V_low
+ 2.148000000e-07 V_low
+ 2.148010000e-07 V_low
+ 2.149000000e-07 V_low
+ 2.149010000e-07 V_hig
+ 2.150000000e-07 V_hig
+ 2.150010000e-07 V_hig
+ 2.151000000e-07 V_hig
+ 2.151010000e-07 V_hig
+ 2.152000000e-07 V_hig
+ 2.152010000e-07 V_hig
+ 2.153000000e-07 V_hig
+ 2.153010000e-07 V_hig
+ 2.154000000e-07 V_hig
+ 2.154010000e-07 V_hig
+ 2.155000000e-07 V_hig
+ 2.155010000e-07 V_hig
+ 2.156000000e-07 V_hig
+ 2.156010000e-07 V_hig
+ 2.157000000e-07 V_hig
+ 2.157010000e-07 V_hig
+ 2.158000000e-07 V_hig
+ 2.158010000e-07 V_hig
+ 2.159000000e-07 V_hig
+ 2.159010000e-07 V_low
+ 2.160000000e-07 V_low
+ 2.160010000e-07 V_low
+ 2.161000000e-07 V_low
+ 2.161010000e-07 V_low
+ 2.162000000e-07 V_low
+ 2.162010000e-07 V_low
+ 2.163000000e-07 V_low
+ 2.163010000e-07 V_low
+ 2.164000000e-07 V_low
+ 2.164010000e-07 V_low
+ 2.165000000e-07 V_low
+ 2.165010000e-07 V_low
+ 2.166000000e-07 V_low
+ 2.166010000e-07 V_low
+ 2.167000000e-07 V_low
+ 2.167010000e-07 V_low
+ 2.168000000e-07 V_low
+ 2.168010000e-07 V_low
+ 2.169000000e-07 V_low
+ 2.169010000e-07 V_low
+ 2.170000000e-07 V_low
+ 2.170010000e-07 V_low
+ 2.171000000e-07 V_low
+ 2.171010000e-07 V_low
+ 2.172000000e-07 V_low
+ 2.172010000e-07 V_low
+ 2.173000000e-07 V_low
+ 2.173010000e-07 V_low
+ 2.174000000e-07 V_low
+ 2.174010000e-07 V_low
+ 2.175000000e-07 V_low
+ 2.175010000e-07 V_low
+ 2.176000000e-07 V_low
+ 2.176010000e-07 V_low
+ 2.177000000e-07 V_low
+ 2.177010000e-07 V_low
+ 2.178000000e-07 V_low
+ 2.178010000e-07 V_low
+ 2.179000000e-07 V_low
+ 2.179010000e-07 V_hig
+ 2.180000000e-07 V_hig
+ 2.180010000e-07 V_hig
+ 2.181000000e-07 V_hig
+ 2.181010000e-07 V_hig
+ 2.182000000e-07 V_hig
+ 2.182010000e-07 V_hig
+ 2.183000000e-07 V_hig
+ 2.183010000e-07 V_hig
+ 2.184000000e-07 V_hig
+ 2.184010000e-07 V_hig
+ 2.185000000e-07 V_hig
+ 2.185010000e-07 V_hig
+ 2.186000000e-07 V_hig
+ 2.186010000e-07 V_hig
+ 2.187000000e-07 V_hig
+ 2.187010000e-07 V_hig
+ 2.188000000e-07 V_hig
+ 2.188010000e-07 V_hig
+ 2.189000000e-07 V_hig
+ 2.189010000e-07 V_hig
+ 2.190000000e-07 V_hig
+ 2.190010000e-07 V_hig
+ 2.191000000e-07 V_hig
+ 2.191010000e-07 V_hig
+ 2.192000000e-07 V_hig
+ 2.192010000e-07 V_hig
+ 2.193000000e-07 V_hig
+ 2.193010000e-07 V_hig
+ 2.194000000e-07 V_hig
+ 2.194010000e-07 V_hig
+ 2.195000000e-07 V_hig
+ 2.195010000e-07 V_hig
+ 2.196000000e-07 V_hig
+ 2.196010000e-07 V_hig
+ 2.197000000e-07 V_hig
+ 2.197010000e-07 V_hig
+ 2.198000000e-07 V_hig
+ 2.198010000e-07 V_hig
+ 2.199000000e-07 V_hig
+ 2.199010000e-07 V_hig
+ 2.200000000e-07 V_hig
+ 2.200010000e-07 V_hig
+ 2.201000000e-07 V_hig
+ 2.201010000e-07 V_hig
+ 2.202000000e-07 V_hig
+ 2.202010000e-07 V_hig
+ 2.203000000e-07 V_hig
+ 2.203010000e-07 V_hig
+ 2.204000000e-07 V_hig
+ 2.204010000e-07 V_hig
+ 2.205000000e-07 V_hig
+ 2.205010000e-07 V_hig
+ 2.206000000e-07 V_hig
+ 2.206010000e-07 V_hig
+ 2.207000000e-07 V_hig
+ 2.207010000e-07 V_hig
+ 2.208000000e-07 V_hig
+ 2.208010000e-07 V_hig
+ 2.209000000e-07 V_hig
+ 2.209010000e-07 V_low
+ 2.210000000e-07 V_low
+ 2.210010000e-07 V_low
+ 2.211000000e-07 V_low
+ 2.211010000e-07 V_low
+ 2.212000000e-07 V_low
+ 2.212010000e-07 V_low
+ 2.213000000e-07 V_low
+ 2.213010000e-07 V_low
+ 2.214000000e-07 V_low
+ 2.214010000e-07 V_low
+ 2.215000000e-07 V_low
+ 2.215010000e-07 V_low
+ 2.216000000e-07 V_low
+ 2.216010000e-07 V_low
+ 2.217000000e-07 V_low
+ 2.217010000e-07 V_low
+ 2.218000000e-07 V_low
+ 2.218010000e-07 V_low
+ 2.219000000e-07 V_low
+ 2.219010000e-07 V_low
+ 2.220000000e-07 V_low
+ 2.220010000e-07 V_low
+ 2.221000000e-07 V_low
+ 2.221010000e-07 V_low
+ 2.222000000e-07 V_low
+ 2.222010000e-07 V_low
+ 2.223000000e-07 V_low
+ 2.223010000e-07 V_low
+ 2.224000000e-07 V_low
+ 2.224010000e-07 V_low
+ 2.225000000e-07 V_low
+ 2.225010000e-07 V_low
+ 2.226000000e-07 V_low
+ 2.226010000e-07 V_low
+ 2.227000000e-07 V_low
+ 2.227010000e-07 V_low
+ 2.228000000e-07 V_low
+ 2.228010000e-07 V_low
+ 2.229000000e-07 V_low
+ 2.229010000e-07 V_low
+ 2.230000000e-07 V_low
+ 2.230010000e-07 V_low
+ 2.231000000e-07 V_low
+ 2.231010000e-07 V_low
+ 2.232000000e-07 V_low
+ 2.232010000e-07 V_low
+ 2.233000000e-07 V_low
+ 2.233010000e-07 V_low
+ 2.234000000e-07 V_low
+ 2.234010000e-07 V_low
+ 2.235000000e-07 V_low
+ 2.235010000e-07 V_low
+ 2.236000000e-07 V_low
+ 2.236010000e-07 V_low
+ 2.237000000e-07 V_low
+ 2.237010000e-07 V_low
+ 2.238000000e-07 V_low
+ 2.238010000e-07 V_low
+ 2.239000000e-07 V_low
+ 2.239010000e-07 V_low
+ 2.240000000e-07 V_low
+ 2.240010000e-07 V_low
+ 2.241000000e-07 V_low
+ 2.241010000e-07 V_low
+ 2.242000000e-07 V_low
+ 2.242010000e-07 V_low
+ 2.243000000e-07 V_low
+ 2.243010000e-07 V_low
+ 2.244000000e-07 V_low
+ 2.244010000e-07 V_low
+ 2.245000000e-07 V_low
+ 2.245010000e-07 V_low
+ 2.246000000e-07 V_low
+ 2.246010000e-07 V_low
+ 2.247000000e-07 V_low
+ 2.247010000e-07 V_low
+ 2.248000000e-07 V_low
+ 2.248010000e-07 V_low
+ 2.249000000e-07 V_low
+ 2.249010000e-07 V_hig
+ 2.250000000e-07 V_hig
+ 2.250010000e-07 V_hig
+ 2.251000000e-07 V_hig
+ 2.251010000e-07 V_hig
+ 2.252000000e-07 V_hig
+ 2.252010000e-07 V_hig
+ 2.253000000e-07 V_hig
+ 2.253010000e-07 V_hig
+ 2.254000000e-07 V_hig
+ 2.254010000e-07 V_hig
+ 2.255000000e-07 V_hig
+ 2.255010000e-07 V_hig
+ 2.256000000e-07 V_hig
+ 2.256010000e-07 V_hig
+ 2.257000000e-07 V_hig
+ 2.257010000e-07 V_hig
+ 2.258000000e-07 V_hig
+ 2.258010000e-07 V_hig
+ 2.259000000e-07 V_hig
+ 2.259010000e-07 V_low
+ 2.260000000e-07 V_low
+ 2.260010000e-07 V_low
+ 2.261000000e-07 V_low
+ 2.261010000e-07 V_low
+ 2.262000000e-07 V_low
+ 2.262010000e-07 V_low
+ 2.263000000e-07 V_low
+ 2.263010000e-07 V_low
+ 2.264000000e-07 V_low
+ 2.264010000e-07 V_low
+ 2.265000000e-07 V_low
+ 2.265010000e-07 V_low
+ 2.266000000e-07 V_low
+ 2.266010000e-07 V_low
+ 2.267000000e-07 V_low
+ 2.267010000e-07 V_low
+ 2.268000000e-07 V_low
+ 2.268010000e-07 V_low
+ 2.269000000e-07 V_low
+ 2.269010000e-07 V_low
+ 2.270000000e-07 V_low
+ 2.270010000e-07 V_low
+ 2.271000000e-07 V_low
+ 2.271010000e-07 V_low
+ 2.272000000e-07 V_low
+ 2.272010000e-07 V_low
+ 2.273000000e-07 V_low
+ 2.273010000e-07 V_low
+ 2.274000000e-07 V_low
+ 2.274010000e-07 V_low
+ 2.275000000e-07 V_low
+ 2.275010000e-07 V_low
+ 2.276000000e-07 V_low
+ 2.276010000e-07 V_low
+ 2.277000000e-07 V_low
+ 2.277010000e-07 V_low
+ 2.278000000e-07 V_low
+ 2.278010000e-07 V_low
+ 2.279000000e-07 V_low
+ 2.279010000e-07 V_hig
+ 2.280000000e-07 V_hig
+ 2.280010000e-07 V_hig
+ 2.281000000e-07 V_hig
+ 2.281010000e-07 V_hig
+ 2.282000000e-07 V_hig
+ 2.282010000e-07 V_hig
+ 2.283000000e-07 V_hig
+ 2.283010000e-07 V_hig
+ 2.284000000e-07 V_hig
+ 2.284010000e-07 V_hig
+ 2.285000000e-07 V_hig
+ 2.285010000e-07 V_hig
+ 2.286000000e-07 V_hig
+ 2.286010000e-07 V_hig
+ 2.287000000e-07 V_hig
+ 2.287010000e-07 V_hig
+ 2.288000000e-07 V_hig
+ 2.288010000e-07 V_hig
+ 2.289000000e-07 V_hig
+ 2.289010000e-07 V_hig
+ 2.290000000e-07 V_hig
+ 2.290010000e-07 V_hig
+ 2.291000000e-07 V_hig
+ 2.291010000e-07 V_hig
+ 2.292000000e-07 V_hig
+ 2.292010000e-07 V_hig
+ 2.293000000e-07 V_hig
+ 2.293010000e-07 V_hig
+ 2.294000000e-07 V_hig
+ 2.294010000e-07 V_hig
+ 2.295000000e-07 V_hig
+ 2.295010000e-07 V_hig
+ 2.296000000e-07 V_hig
+ 2.296010000e-07 V_hig
+ 2.297000000e-07 V_hig
+ 2.297010000e-07 V_hig
+ 2.298000000e-07 V_hig
+ 2.298010000e-07 V_hig
+ 2.299000000e-07 V_hig
+ 2.299010000e-07 V_low
+ 2.300000000e-07 V_low
+ 2.300010000e-07 V_low
+ 2.301000000e-07 V_low
+ 2.301010000e-07 V_low
+ 2.302000000e-07 V_low
+ 2.302010000e-07 V_low
+ 2.303000000e-07 V_low
+ 2.303010000e-07 V_low
+ 2.304000000e-07 V_low
+ 2.304010000e-07 V_low
+ 2.305000000e-07 V_low
+ 2.305010000e-07 V_low
+ 2.306000000e-07 V_low
+ 2.306010000e-07 V_low
+ 2.307000000e-07 V_low
+ 2.307010000e-07 V_low
+ 2.308000000e-07 V_low
+ 2.308010000e-07 V_low
+ 2.309000000e-07 V_low
+ 2.309010000e-07 V_hig
+ 2.310000000e-07 V_hig
+ 2.310010000e-07 V_hig
+ 2.311000000e-07 V_hig
+ 2.311010000e-07 V_hig
+ 2.312000000e-07 V_hig
+ 2.312010000e-07 V_hig
+ 2.313000000e-07 V_hig
+ 2.313010000e-07 V_hig
+ 2.314000000e-07 V_hig
+ 2.314010000e-07 V_hig
+ 2.315000000e-07 V_hig
+ 2.315010000e-07 V_hig
+ 2.316000000e-07 V_hig
+ 2.316010000e-07 V_hig
+ 2.317000000e-07 V_hig
+ 2.317010000e-07 V_hig
+ 2.318000000e-07 V_hig
+ 2.318010000e-07 V_hig
+ 2.319000000e-07 V_hig
+ 2.319010000e-07 V_hig
+ 2.320000000e-07 V_hig
+ 2.320010000e-07 V_hig
+ 2.321000000e-07 V_hig
+ 2.321010000e-07 V_hig
+ 2.322000000e-07 V_hig
+ 2.322010000e-07 V_hig
+ 2.323000000e-07 V_hig
+ 2.323010000e-07 V_hig
+ 2.324000000e-07 V_hig
+ 2.324010000e-07 V_hig
+ 2.325000000e-07 V_hig
+ 2.325010000e-07 V_hig
+ 2.326000000e-07 V_hig
+ 2.326010000e-07 V_hig
+ 2.327000000e-07 V_hig
+ 2.327010000e-07 V_hig
+ 2.328000000e-07 V_hig
+ 2.328010000e-07 V_hig
+ 2.329000000e-07 V_hig
+ 2.329010000e-07 V_low
+ 2.330000000e-07 V_low
+ 2.330010000e-07 V_low
+ 2.331000000e-07 V_low
+ 2.331010000e-07 V_low
+ 2.332000000e-07 V_low
+ 2.332010000e-07 V_low
+ 2.333000000e-07 V_low
+ 2.333010000e-07 V_low
+ 2.334000000e-07 V_low
+ 2.334010000e-07 V_low
+ 2.335000000e-07 V_low
+ 2.335010000e-07 V_low
+ 2.336000000e-07 V_low
+ 2.336010000e-07 V_low
+ 2.337000000e-07 V_low
+ 2.337010000e-07 V_low
+ 2.338000000e-07 V_low
+ 2.338010000e-07 V_low
+ 2.339000000e-07 V_low
+ 2.339010000e-07 V_low
+ 2.340000000e-07 V_low
+ 2.340010000e-07 V_low
+ 2.341000000e-07 V_low
+ 2.341010000e-07 V_low
+ 2.342000000e-07 V_low
+ 2.342010000e-07 V_low
+ 2.343000000e-07 V_low
+ 2.343010000e-07 V_low
+ 2.344000000e-07 V_low
+ 2.344010000e-07 V_low
+ 2.345000000e-07 V_low
+ 2.345010000e-07 V_low
+ 2.346000000e-07 V_low
+ 2.346010000e-07 V_low
+ 2.347000000e-07 V_low
+ 2.347010000e-07 V_low
+ 2.348000000e-07 V_low
+ 2.348010000e-07 V_low
+ 2.349000000e-07 V_low
+ 2.349010000e-07 V_low
+ 2.350000000e-07 V_low
+ 2.350010000e-07 V_low
+ 2.351000000e-07 V_low
+ 2.351010000e-07 V_low
+ 2.352000000e-07 V_low
+ 2.352010000e-07 V_low
+ 2.353000000e-07 V_low
+ 2.353010000e-07 V_low
+ 2.354000000e-07 V_low
+ 2.354010000e-07 V_low
+ 2.355000000e-07 V_low
+ 2.355010000e-07 V_low
+ 2.356000000e-07 V_low
+ 2.356010000e-07 V_low
+ 2.357000000e-07 V_low
+ 2.357010000e-07 V_low
+ 2.358000000e-07 V_low
+ 2.358010000e-07 V_low
+ 2.359000000e-07 V_low
+ 2.359010000e-07 V_low
+ 2.360000000e-07 V_low
+ 2.360010000e-07 V_low
+ 2.361000000e-07 V_low
+ 2.361010000e-07 V_low
+ 2.362000000e-07 V_low
+ 2.362010000e-07 V_low
+ 2.363000000e-07 V_low
+ 2.363010000e-07 V_low
+ 2.364000000e-07 V_low
+ 2.364010000e-07 V_low
+ 2.365000000e-07 V_low
+ 2.365010000e-07 V_low
+ 2.366000000e-07 V_low
+ 2.366010000e-07 V_low
+ 2.367000000e-07 V_low
+ 2.367010000e-07 V_low
+ 2.368000000e-07 V_low
+ 2.368010000e-07 V_low
+ 2.369000000e-07 V_low
+ 2.369010000e-07 V_hig
+ 2.370000000e-07 V_hig
+ 2.370010000e-07 V_hig
+ 2.371000000e-07 V_hig
+ 2.371010000e-07 V_hig
+ 2.372000000e-07 V_hig
+ 2.372010000e-07 V_hig
+ 2.373000000e-07 V_hig
+ 2.373010000e-07 V_hig
+ 2.374000000e-07 V_hig
+ 2.374010000e-07 V_hig
+ 2.375000000e-07 V_hig
+ 2.375010000e-07 V_hig
+ 2.376000000e-07 V_hig
+ 2.376010000e-07 V_hig
+ 2.377000000e-07 V_hig
+ 2.377010000e-07 V_hig
+ 2.378000000e-07 V_hig
+ 2.378010000e-07 V_hig
+ 2.379000000e-07 V_hig
+ 2.379010000e-07 V_low
+ 2.380000000e-07 V_low
+ 2.380010000e-07 V_low
+ 2.381000000e-07 V_low
+ 2.381010000e-07 V_low
+ 2.382000000e-07 V_low
+ 2.382010000e-07 V_low
+ 2.383000000e-07 V_low
+ 2.383010000e-07 V_low
+ 2.384000000e-07 V_low
+ 2.384010000e-07 V_low
+ 2.385000000e-07 V_low
+ 2.385010000e-07 V_low
+ 2.386000000e-07 V_low
+ 2.386010000e-07 V_low
+ 2.387000000e-07 V_low
+ 2.387010000e-07 V_low
+ 2.388000000e-07 V_low
+ 2.388010000e-07 V_low
+ 2.389000000e-07 V_low
+ 2.389010000e-07 V_hig
+ 2.390000000e-07 V_hig
+ 2.390010000e-07 V_hig
+ 2.391000000e-07 V_hig
+ 2.391010000e-07 V_hig
+ 2.392000000e-07 V_hig
+ 2.392010000e-07 V_hig
+ 2.393000000e-07 V_hig
+ 2.393010000e-07 V_hig
+ 2.394000000e-07 V_hig
+ 2.394010000e-07 V_hig
+ 2.395000000e-07 V_hig
+ 2.395010000e-07 V_hig
+ 2.396000000e-07 V_hig
+ 2.396010000e-07 V_hig
+ 2.397000000e-07 V_hig
+ 2.397010000e-07 V_hig
+ 2.398000000e-07 V_hig
+ 2.398010000e-07 V_hig
+ 2.399000000e-07 V_hig
+ 2.399010000e-07 V_low
+ 2.400000000e-07 V_low
+ 2.400010000e-07 V_low
+ 2.401000000e-07 V_low
+ 2.401010000e-07 V_low
+ 2.402000000e-07 V_low
+ 2.402010000e-07 V_low
+ 2.403000000e-07 V_low
+ 2.403010000e-07 V_low
+ 2.404000000e-07 V_low
+ 2.404010000e-07 V_low
+ 2.405000000e-07 V_low
+ 2.405010000e-07 V_low
+ 2.406000000e-07 V_low
+ 2.406010000e-07 V_low
+ 2.407000000e-07 V_low
+ 2.407010000e-07 V_low
+ 2.408000000e-07 V_low
+ 2.408010000e-07 V_low
+ 2.409000000e-07 V_low
+ 2.409010000e-07 V_low
+ 2.410000000e-07 V_low
+ 2.410010000e-07 V_low
+ 2.411000000e-07 V_low
+ 2.411010000e-07 V_low
+ 2.412000000e-07 V_low
+ 2.412010000e-07 V_low
+ 2.413000000e-07 V_low
+ 2.413010000e-07 V_low
+ 2.414000000e-07 V_low
+ 2.414010000e-07 V_low
+ 2.415000000e-07 V_low
+ 2.415010000e-07 V_low
+ 2.416000000e-07 V_low
+ 2.416010000e-07 V_low
+ 2.417000000e-07 V_low
+ 2.417010000e-07 V_low
+ 2.418000000e-07 V_low
+ 2.418010000e-07 V_low
+ 2.419000000e-07 V_low
+ 2.419010000e-07 V_low
+ 2.420000000e-07 V_low
+ 2.420010000e-07 V_low
+ 2.421000000e-07 V_low
+ 2.421010000e-07 V_low
+ 2.422000000e-07 V_low
+ 2.422010000e-07 V_low
+ 2.423000000e-07 V_low
+ 2.423010000e-07 V_low
+ 2.424000000e-07 V_low
+ 2.424010000e-07 V_low
+ 2.425000000e-07 V_low
+ 2.425010000e-07 V_low
+ 2.426000000e-07 V_low
+ 2.426010000e-07 V_low
+ 2.427000000e-07 V_low
+ 2.427010000e-07 V_low
+ 2.428000000e-07 V_low
+ 2.428010000e-07 V_low
+ 2.429000000e-07 V_low
+ 2.429010000e-07 V_low
+ 2.430000000e-07 V_low
+ 2.430010000e-07 V_low
+ 2.431000000e-07 V_low
+ 2.431010000e-07 V_low
+ 2.432000000e-07 V_low
+ 2.432010000e-07 V_low
+ 2.433000000e-07 V_low
+ 2.433010000e-07 V_low
+ 2.434000000e-07 V_low
+ 2.434010000e-07 V_low
+ 2.435000000e-07 V_low
+ 2.435010000e-07 V_low
+ 2.436000000e-07 V_low
+ 2.436010000e-07 V_low
+ 2.437000000e-07 V_low
+ 2.437010000e-07 V_low
+ 2.438000000e-07 V_low
+ 2.438010000e-07 V_low
+ 2.439000000e-07 V_low
+ 2.439010000e-07 V_hig
+ 2.440000000e-07 V_hig
+ 2.440010000e-07 V_hig
+ 2.441000000e-07 V_hig
+ 2.441010000e-07 V_hig
+ 2.442000000e-07 V_hig
+ 2.442010000e-07 V_hig
+ 2.443000000e-07 V_hig
+ 2.443010000e-07 V_hig
+ 2.444000000e-07 V_hig
+ 2.444010000e-07 V_hig
+ 2.445000000e-07 V_hig
+ 2.445010000e-07 V_hig
+ 2.446000000e-07 V_hig
+ 2.446010000e-07 V_hig
+ 2.447000000e-07 V_hig
+ 2.447010000e-07 V_hig
+ 2.448000000e-07 V_hig
+ 2.448010000e-07 V_hig
+ 2.449000000e-07 V_hig
+ 2.449010000e-07 V_low
+ 2.450000000e-07 V_low
+ 2.450010000e-07 V_low
+ 2.451000000e-07 V_low
+ 2.451010000e-07 V_low
+ 2.452000000e-07 V_low
+ 2.452010000e-07 V_low
+ 2.453000000e-07 V_low
+ 2.453010000e-07 V_low
+ 2.454000000e-07 V_low
+ 2.454010000e-07 V_low
+ 2.455000000e-07 V_low
+ 2.455010000e-07 V_low
+ 2.456000000e-07 V_low
+ 2.456010000e-07 V_low
+ 2.457000000e-07 V_low
+ 2.457010000e-07 V_low
+ 2.458000000e-07 V_low
+ 2.458010000e-07 V_low
+ 2.459000000e-07 V_low
+ 2.459010000e-07 V_low
+ 2.460000000e-07 V_low
+ 2.460010000e-07 V_low
+ 2.461000000e-07 V_low
+ 2.461010000e-07 V_low
+ 2.462000000e-07 V_low
+ 2.462010000e-07 V_low
+ 2.463000000e-07 V_low
+ 2.463010000e-07 V_low
+ 2.464000000e-07 V_low
+ 2.464010000e-07 V_low
+ 2.465000000e-07 V_low
+ 2.465010000e-07 V_low
+ 2.466000000e-07 V_low
+ 2.466010000e-07 V_low
+ 2.467000000e-07 V_low
+ 2.467010000e-07 V_low
+ 2.468000000e-07 V_low
+ 2.468010000e-07 V_low
+ 2.469000000e-07 V_low
+ 2.469010000e-07 V_low
+ 2.470000000e-07 V_low
+ 2.470010000e-07 V_low
+ 2.471000000e-07 V_low
+ 2.471010000e-07 V_low
+ 2.472000000e-07 V_low
+ 2.472010000e-07 V_low
+ 2.473000000e-07 V_low
+ 2.473010000e-07 V_low
+ 2.474000000e-07 V_low
+ 2.474010000e-07 V_low
+ 2.475000000e-07 V_low
+ 2.475010000e-07 V_low
+ 2.476000000e-07 V_low
+ 2.476010000e-07 V_low
+ 2.477000000e-07 V_low
+ 2.477010000e-07 V_low
+ 2.478000000e-07 V_low
+ 2.478010000e-07 V_low
+ 2.479000000e-07 V_low
+ 2.479010000e-07 V_low
+ 2.480000000e-07 V_low
+ 2.480010000e-07 V_low
+ 2.481000000e-07 V_low
+ 2.481010000e-07 V_low
+ 2.482000000e-07 V_low
+ 2.482010000e-07 V_low
+ 2.483000000e-07 V_low
+ 2.483010000e-07 V_low
+ 2.484000000e-07 V_low
+ 2.484010000e-07 V_low
+ 2.485000000e-07 V_low
+ 2.485010000e-07 V_low
+ 2.486000000e-07 V_low
+ 2.486010000e-07 V_low
+ 2.487000000e-07 V_low
+ 2.487010000e-07 V_low
+ 2.488000000e-07 V_low
+ 2.488010000e-07 V_low
+ 2.489000000e-07 V_low
+ 2.489010000e-07 V_hig
+ 2.490000000e-07 V_hig
+ 2.490010000e-07 V_hig
+ 2.491000000e-07 V_hig
+ 2.491010000e-07 V_hig
+ 2.492000000e-07 V_hig
+ 2.492010000e-07 V_hig
+ 2.493000000e-07 V_hig
+ 2.493010000e-07 V_hig
+ 2.494000000e-07 V_hig
+ 2.494010000e-07 V_hig
+ 2.495000000e-07 V_hig
+ 2.495010000e-07 V_hig
+ 2.496000000e-07 V_hig
+ 2.496010000e-07 V_hig
+ 2.497000000e-07 V_hig
+ 2.497010000e-07 V_hig
+ 2.498000000e-07 V_hig
+ 2.498010000e-07 V_hig
+ 2.499000000e-07 V_hig
+ 2.499010000e-07 V_hig
+ 2.500000000e-07 V_hig
+ 2.500010000e-07 V_hig
+ 2.501000000e-07 V_hig
+ 2.501010000e-07 V_hig
+ 2.502000000e-07 V_hig
+ 2.502010000e-07 V_hig
+ 2.503000000e-07 V_hig
+ 2.503010000e-07 V_hig
+ 2.504000000e-07 V_hig
+ 2.504010000e-07 V_hig
+ 2.505000000e-07 V_hig
+ 2.505010000e-07 V_hig
+ 2.506000000e-07 V_hig
+ 2.506010000e-07 V_hig
+ 2.507000000e-07 V_hig
+ 2.507010000e-07 V_hig
+ 2.508000000e-07 V_hig
+ 2.508010000e-07 V_hig
+ 2.509000000e-07 V_hig
+ 2.509010000e-07 V_low
+ 2.510000000e-07 V_low
+ 2.510010000e-07 V_low
+ 2.511000000e-07 V_low
+ 2.511010000e-07 V_low
+ 2.512000000e-07 V_low
+ 2.512010000e-07 V_low
+ 2.513000000e-07 V_low
+ 2.513010000e-07 V_low
+ 2.514000000e-07 V_low
+ 2.514010000e-07 V_low
+ 2.515000000e-07 V_low
+ 2.515010000e-07 V_low
+ 2.516000000e-07 V_low
+ 2.516010000e-07 V_low
+ 2.517000000e-07 V_low
+ 2.517010000e-07 V_low
+ 2.518000000e-07 V_low
+ 2.518010000e-07 V_low
+ 2.519000000e-07 V_low
+ 2.519010000e-07 V_low
+ 2.520000000e-07 V_low
+ 2.520010000e-07 V_low
+ 2.521000000e-07 V_low
+ 2.521010000e-07 V_low
+ 2.522000000e-07 V_low
+ 2.522010000e-07 V_low
+ 2.523000000e-07 V_low
+ 2.523010000e-07 V_low
+ 2.524000000e-07 V_low
+ 2.524010000e-07 V_low
+ 2.525000000e-07 V_low
+ 2.525010000e-07 V_low
+ 2.526000000e-07 V_low
+ 2.526010000e-07 V_low
+ 2.527000000e-07 V_low
+ 2.527010000e-07 V_low
+ 2.528000000e-07 V_low
+ 2.528010000e-07 V_low
+ 2.529000000e-07 V_low
+ 2.529010000e-07 V_low
+ 2.530000000e-07 V_low
+ 2.530010000e-07 V_low
+ 2.531000000e-07 V_low
+ 2.531010000e-07 V_low
+ 2.532000000e-07 V_low
+ 2.532010000e-07 V_low
+ 2.533000000e-07 V_low
+ 2.533010000e-07 V_low
+ 2.534000000e-07 V_low
+ 2.534010000e-07 V_low
+ 2.535000000e-07 V_low
+ 2.535010000e-07 V_low
+ 2.536000000e-07 V_low
+ 2.536010000e-07 V_low
+ 2.537000000e-07 V_low
+ 2.537010000e-07 V_low
+ 2.538000000e-07 V_low
+ 2.538010000e-07 V_low
+ 2.539000000e-07 V_low
+ 2.539010000e-07 V_low
+ 2.540000000e-07 V_low
+ 2.540010000e-07 V_low
+ 2.541000000e-07 V_low
+ 2.541010000e-07 V_low
+ 2.542000000e-07 V_low
+ 2.542010000e-07 V_low
+ 2.543000000e-07 V_low
+ 2.543010000e-07 V_low
+ 2.544000000e-07 V_low
+ 2.544010000e-07 V_low
+ 2.545000000e-07 V_low
+ 2.545010000e-07 V_low
+ 2.546000000e-07 V_low
+ 2.546010000e-07 V_low
+ 2.547000000e-07 V_low
+ 2.547010000e-07 V_low
+ 2.548000000e-07 V_low
+ 2.548010000e-07 V_low
+ 2.549000000e-07 V_low
+ 2.549010000e-07 V_hig
+ 2.550000000e-07 V_hig
+ 2.550010000e-07 V_hig
+ 2.551000000e-07 V_hig
+ 2.551010000e-07 V_hig
+ 2.552000000e-07 V_hig
+ 2.552010000e-07 V_hig
+ 2.553000000e-07 V_hig
+ 2.553010000e-07 V_hig
+ 2.554000000e-07 V_hig
+ 2.554010000e-07 V_hig
+ 2.555000000e-07 V_hig
+ 2.555010000e-07 V_hig
+ 2.556000000e-07 V_hig
+ 2.556010000e-07 V_hig
+ 2.557000000e-07 V_hig
+ 2.557010000e-07 V_hig
+ 2.558000000e-07 V_hig
+ 2.558010000e-07 V_hig
+ 2.559000000e-07 V_hig
+ 2.559010000e-07 V_low
+ 2.560000000e-07 V_low
+ 2.560010000e-07 V_low
+ 2.561000000e-07 V_low
+ 2.561010000e-07 V_low
+ 2.562000000e-07 V_low
+ 2.562010000e-07 V_low
+ 2.563000000e-07 V_low
+ 2.563010000e-07 V_low
+ 2.564000000e-07 V_low
+ 2.564010000e-07 V_low
+ 2.565000000e-07 V_low
+ 2.565010000e-07 V_low
+ 2.566000000e-07 V_low
+ 2.566010000e-07 V_low
+ 2.567000000e-07 V_low
+ 2.567010000e-07 V_low
+ 2.568000000e-07 V_low
+ 2.568010000e-07 V_low
+ 2.569000000e-07 V_low
+ 2.569010000e-07 V_hig
+ 2.570000000e-07 V_hig
+ 2.570010000e-07 V_hig
+ 2.571000000e-07 V_hig
+ 2.571010000e-07 V_hig
+ 2.572000000e-07 V_hig
+ 2.572010000e-07 V_hig
+ 2.573000000e-07 V_hig
+ 2.573010000e-07 V_hig
+ 2.574000000e-07 V_hig
+ 2.574010000e-07 V_hig
+ 2.575000000e-07 V_hig
+ 2.575010000e-07 V_hig
+ 2.576000000e-07 V_hig
+ 2.576010000e-07 V_hig
+ 2.577000000e-07 V_hig
+ 2.577010000e-07 V_hig
+ 2.578000000e-07 V_hig
+ 2.578010000e-07 V_hig
+ 2.579000000e-07 V_hig
+ 2.579010000e-07 V_low
+ 2.580000000e-07 V_low
+ 2.580010000e-07 V_low
+ 2.581000000e-07 V_low
+ 2.581010000e-07 V_low
+ 2.582000000e-07 V_low
+ 2.582010000e-07 V_low
+ 2.583000000e-07 V_low
+ 2.583010000e-07 V_low
+ 2.584000000e-07 V_low
+ 2.584010000e-07 V_low
+ 2.585000000e-07 V_low
+ 2.585010000e-07 V_low
+ 2.586000000e-07 V_low
+ 2.586010000e-07 V_low
+ 2.587000000e-07 V_low
+ 2.587010000e-07 V_low
+ 2.588000000e-07 V_low
+ 2.588010000e-07 V_low
+ 2.589000000e-07 V_low
+ 2.589010000e-07 V_hig
+ 2.590000000e-07 V_hig
+ 2.590010000e-07 V_hig
+ 2.591000000e-07 V_hig
+ 2.591010000e-07 V_hig
+ 2.592000000e-07 V_hig
+ 2.592010000e-07 V_hig
+ 2.593000000e-07 V_hig
+ 2.593010000e-07 V_hig
+ 2.594000000e-07 V_hig
+ 2.594010000e-07 V_hig
+ 2.595000000e-07 V_hig
+ 2.595010000e-07 V_hig
+ 2.596000000e-07 V_hig
+ 2.596010000e-07 V_hig
+ 2.597000000e-07 V_hig
+ 2.597010000e-07 V_hig
+ 2.598000000e-07 V_hig
+ 2.598010000e-07 V_hig
+ 2.599000000e-07 V_hig
+ 2.599010000e-07 V_hig
+ 2.600000000e-07 V_hig
+ 2.600010000e-07 V_hig
+ 2.601000000e-07 V_hig
+ 2.601010000e-07 V_hig
+ 2.602000000e-07 V_hig
+ 2.602010000e-07 V_hig
+ 2.603000000e-07 V_hig
+ 2.603010000e-07 V_hig
+ 2.604000000e-07 V_hig
+ 2.604010000e-07 V_hig
+ 2.605000000e-07 V_hig
+ 2.605010000e-07 V_hig
+ 2.606000000e-07 V_hig
+ 2.606010000e-07 V_hig
+ 2.607000000e-07 V_hig
+ 2.607010000e-07 V_hig
+ 2.608000000e-07 V_hig
+ 2.608010000e-07 V_hig
+ 2.609000000e-07 V_hig
+ 2.609010000e-07 V_hig
+ 2.610000000e-07 V_hig
+ 2.610010000e-07 V_hig
+ 2.611000000e-07 V_hig
+ 2.611010000e-07 V_hig
+ 2.612000000e-07 V_hig
+ 2.612010000e-07 V_hig
+ 2.613000000e-07 V_hig
+ 2.613010000e-07 V_hig
+ 2.614000000e-07 V_hig
+ 2.614010000e-07 V_hig
+ 2.615000000e-07 V_hig
+ 2.615010000e-07 V_hig
+ 2.616000000e-07 V_hig
+ 2.616010000e-07 V_hig
+ 2.617000000e-07 V_hig
+ 2.617010000e-07 V_hig
+ 2.618000000e-07 V_hig
+ 2.618010000e-07 V_hig
+ 2.619000000e-07 V_hig
+ 2.619010000e-07 V_hig
+ 2.620000000e-07 V_hig
+ 2.620010000e-07 V_hig
+ 2.621000000e-07 V_hig
+ 2.621010000e-07 V_hig
+ 2.622000000e-07 V_hig
+ 2.622010000e-07 V_hig
+ 2.623000000e-07 V_hig
+ 2.623010000e-07 V_hig
+ 2.624000000e-07 V_hig
+ 2.624010000e-07 V_hig
+ 2.625000000e-07 V_hig
+ 2.625010000e-07 V_hig
+ 2.626000000e-07 V_hig
+ 2.626010000e-07 V_hig
+ 2.627000000e-07 V_hig
+ 2.627010000e-07 V_hig
+ 2.628000000e-07 V_hig
+ 2.628010000e-07 V_hig
+ 2.629000000e-07 V_hig
+ 2.629010000e-07 V_hig
+ 2.630000000e-07 V_hig
+ 2.630010000e-07 V_hig
+ 2.631000000e-07 V_hig
+ 2.631010000e-07 V_hig
+ 2.632000000e-07 V_hig
+ 2.632010000e-07 V_hig
+ 2.633000000e-07 V_hig
+ 2.633010000e-07 V_hig
+ 2.634000000e-07 V_hig
+ 2.634010000e-07 V_hig
+ 2.635000000e-07 V_hig
+ 2.635010000e-07 V_hig
+ 2.636000000e-07 V_hig
+ 2.636010000e-07 V_hig
+ 2.637000000e-07 V_hig
+ 2.637010000e-07 V_hig
+ 2.638000000e-07 V_hig
+ 2.638010000e-07 V_hig
+ 2.639000000e-07 V_hig
+ 2.639010000e-07 V_hig
+ 2.640000000e-07 V_hig
+ 2.640010000e-07 V_hig
+ 2.641000000e-07 V_hig
+ 2.641010000e-07 V_hig
+ 2.642000000e-07 V_hig
+ 2.642010000e-07 V_hig
+ 2.643000000e-07 V_hig
+ 2.643010000e-07 V_hig
+ 2.644000000e-07 V_hig
+ 2.644010000e-07 V_hig
+ 2.645000000e-07 V_hig
+ 2.645010000e-07 V_hig
+ 2.646000000e-07 V_hig
+ 2.646010000e-07 V_hig
+ 2.647000000e-07 V_hig
+ 2.647010000e-07 V_hig
+ 2.648000000e-07 V_hig
+ 2.648010000e-07 V_hig
+ 2.649000000e-07 V_hig
+ 2.649010000e-07 V_hig
+ 2.650000000e-07 V_hig
+ 2.650010000e-07 V_hig
+ 2.651000000e-07 V_hig
+ 2.651010000e-07 V_hig
+ 2.652000000e-07 V_hig
+ 2.652010000e-07 V_hig
+ 2.653000000e-07 V_hig
+ 2.653010000e-07 V_hig
+ 2.654000000e-07 V_hig
+ 2.654010000e-07 V_hig
+ 2.655000000e-07 V_hig
+ 2.655010000e-07 V_hig
+ 2.656000000e-07 V_hig
+ 2.656010000e-07 V_hig
+ 2.657000000e-07 V_hig
+ 2.657010000e-07 V_hig
+ 2.658000000e-07 V_hig
+ 2.658010000e-07 V_hig
+ 2.659000000e-07 V_hig
+ 2.659010000e-07 V_low
+ 2.660000000e-07 V_low
+ 2.660010000e-07 V_low
+ 2.661000000e-07 V_low
+ 2.661010000e-07 V_low
+ 2.662000000e-07 V_low
+ 2.662010000e-07 V_low
+ 2.663000000e-07 V_low
+ 2.663010000e-07 V_low
+ 2.664000000e-07 V_low
+ 2.664010000e-07 V_low
+ 2.665000000e-07 V_low
+ 2.665010000e-07 V_low
+ 2.666000000e-07 V_low
+ 2.666010000e-07 V_low
+ 2.667000000e-07 V_low
+ 2.667010000e-07 V_low
+ 2.668000000e-07 V_low
+ 2.668010000e-07 V_low
+ 2.669000000e-07 V_low
+ 2.669010000e-07 V_low
+ 2.670000000e-07 V_low
+ 2.670010000e-07 V_low
+ 2.671000000e-07 V_low
+ 2.671010000e-07 V_low
+ 2.672000000e-07 V_low
+ 2.672010000e-07 V_low
+ 2.673000000e-07 V_low
+ 2.673010000e-07 V_low
+ 2.674000000e-07 V_low
+ 2.674010000e-07 V_low
+ 2.675000000e-07 V_low
+ 2.675010000e-07 V_low
+ 2.676000000e-07 V_low
+ 2.676010000e-07 V_low
+ 2.677000000e-07 V_low
+ 2.677010000e-07 V_low
+ 2.678000000e-07 V_low
+ 2.678010000e-07 V_low
+ 2.679000000e-07 V_low
+ 2.679010000e-07 V_low
+ 2.680000000e-07 V_low
+ 2.680010000e-07 V_low
+ 2.681000000e-07 V_low
+ 2.681010000e-07 V_low
+ 2.682000000e-07 V_low
+ 2.682010000e-07 V_low
+ 2.683000000e-07 V_low
+ 2.683010000e-07 V_low
+ 2.684000000e-07 V_low
+ 2.684010000e-07 V_low
+ 2.685000000e-07 V_low
+ 2.685010000e-07 V_low
+ 2.686000000e-07 V_low
+ 2.686010000e-07 V_low
+ 2.687000000e-07 V_low
+ 2.687010000e-07 V_low
+ 2.688000000e-07 V_low
+ 2.688010000e-07 V_low
+ 2.689000000e-07 V_low
+ 2.689010000e-07 V_low
+ 2.690000000e-07 V_low
+ 2.690010000e-07 V_low
+ 2.691000000e-07 V_low
+ 2.691010000e-07 V_low
+ 2.692000000e-07 V_low
+ 2.692010000e-07 V_low
+ 2.693000000e-07 V_low
+ 2.693010000e-07 V_low
+ 2.694000000e-07 V_low
+ 2.694010000e-07 V_low
+ 2.695000000e-07 V_low
+ 2.695010000e-07 V_low
+ 2.696000000e-07 V_low
+ 2.696010000e-07 V_low
+ 2.697000000e-07 V_low
+ 2.697010000e-07 V_low
+ 2.698000000e-07 V_low
+ 2.698010000e-07 V_low
+ 2.699000000e-07 V_low
+ 2.699010000e-07 V_low
+ 2.700000000e-07 V_low
+ 2.700010000e-07 V_low
+ 2.701000000e-07 V_low
+ 2.701010000e-07 V_low
+ 2.702000000e-07 V_low
+ 2.702010000e-07 V_low
+ 2.703000000e-07 V_low
+ 2.703010000e-07 V_low
+ 2.704000000e-07 V_low
+ 2.704010000e-07 V_low
+ 2.705000000e-07 V_low
+ 2.705010000e-07 V_low
+ 2.706000000e-07 V_low
+ 2.706010000e-07 V_low
+ 2.707000000e-07 V_low
+ 2.707010000e-07 V_low
+ 2.708000000e-07 V_low
+ 2.708010000e-07 V_low
+ 2.709000000e-07 V_low
+ 2.709010000e-07 V_low
+ 2.710000000e-07 V_low
+ 2.710010000e-07 V_low
+ 2.711000000e-07 V_low
+ 2.711010000e-07 V_low
+ 2.712000000e-07 V_low
+ 2.712010000e-07 V_low
+ 2.713000000e-07 V_low
+ 2.713010000e-07 V_low
+ 2.714000000e-07 V_low
+ 2.714010000e-07 V_low
+ 2.715000000e-07 V_low
+ 2.715010000e-07 V_low
+ 2.716000000e-07 V_low
+ 2.716010000e-07 V_low
+ 2.717000000e-07 V_low
+ 2.717010000e-07 V_low
+ 2.718000000e-07 V_low
+ 2.718010000e-07 V_low
+ 2.719000000e-07 V_low
+ 2.719010000e-07 V_low
+ 2.720000000e-07 V_low
+ 2.720010000e-07 V_low
+ 2.721000000e-07 V_low
+ 2.721010000e-07 V_low
+ 2.722000000e-07 V_low
+ 2.722010000e-07 V_low
+ 2.723000000e-07 V_low
+ 2.723010000e-07 V_low
+ 2.724000000e-07 V_low
+ 2.724010000e-07 V_low
+ 2.725000000e-07 V_low
+ 2.725010000e-07 V_low
+ 2.726000000e-07 V_low
+ 2.726010000e-07 V_low
+ 2.727000000e-07 V_low
+ 2.727010000e-07 V_low
+ 2.728000000e-07 V_low
+ 2.728010000e-07 V_low
+ 2.729000000e-07 V_low
+ 2.729010000e-07 V_hig
+ 2.730000000e-07 V_hig
+ 2.730010000e-07 V_hig
+ 2.731000000e-07 V_hig
+ 2.731010000e-07 V_hig
+ 2.732000000e-07 V_hig
+ 2.732010000e-07 V_hig
+ 2.733000000e-07 V_hig
+ 2.733010000e-07 V_hig
+ 2.734000000e-07 V_hig
+ 2.734010000e-07 V_hig
+ 2.735000000e-07 V_hig
+ 2.735010000e-07 V_hig
+ 2.736000000e-07 V_hig
+ 2.736010000e-07 V_hig
+ 2.737000000e-07 V_hig
+ 2.737010000e-07 V_hig
+ 2.738000000e-07 V_hig
+ 2.738010000e-07 V_hig
+ 2.739000000e-07 V_hig
+ 2.739010000e-07 V_hig
+ 2.740000000e-07 V_hig
+ 2.740010000e-07 V_hig
+ 2.741000000e-07 V_hig
+ 2.741010000e-07 V_hig
+ 2.742000000e-07 V_hig
+ 2.742010000e-07 V_hig
+ 2.743000000e-07 V_hig
+ 2.743010000e-07 V_hig
+ 2.744000000e-07 V_hig
+ 2.744010000e-07 V_hig
+ 2.745000000e-07 V_hig
+ 2.745010000e-07 V_hig
+ 2.746000000e-07 V_hig
+ 2.746010000e-07 V_hig
+ 2.747000000e-07 V_hig
+ 2.747010000e-07 V_hig
+ 2.748000000e-07 V_hig
+ 2.748010000e-07 V_hig
+ 2.749000000e-07 V_hig
+ 2.749010000e-07 V_hig
+ 2.750000000e-07 V_hig
+ 2.750010000e-07 V_hig
+ 2.751000000e-07 V_hig
+ 2.751010000e-07 V_hig
+ 2.752000000e-07 V_hig
+ 2.752010000e-07 V_hig
+ 2.753000000e-07 V_hig
+ 2.753010000e-07 V_hig
+ 2.754000000e-07 V_hig
+ 2.754010000e-07 V_hig
+ 2.755000000e-07 V_hig
+ 2.755010000e-07 V_hig
+ 2.756000000e-07 V_hig
+ 2.756010000e-07 V_hig
+ 2.757000000e-07 V_hig
+ 2.757010000e-07 V_hig
+ 2.758000000e-07 V_hig
+ 2.758010000e-07 V_hig
+ 2.759000000e-07 V_hig
+ 2.759010000e-07 V_hig
+ 2.760000000e-07 V_hig
+ 2.760010000e-07 V_hig
+ 2.761000000e-07 V_hig
+ 2.761010000e-07 V_hig
+ 2.762000000e-07 V_hig
+ 2.762010000e-07 V_hig
+ 2.763000000e-07 V_hig
+ 2.763010000e-07 V_hig
+ 2.764000000e-07 V_hig
+ 2.764010000e-07 V_hig
+ 2.765000000e-07 V_hig
+ 2.765010000e-07 V_hig
+ 2.766000000e-07 V_hig
+ 2.766010000e-07 V_hig
+ 2.767000000e-07 V_hig
+ 2.767010000e-07 V_hig
+ 2.768000000e-07 V_hig
+ 2.768010000e-07 V_hig
+ 2.769000000e-07 V_hig
+ 2.769010000e-07 V_hig
+ 2.770000000e-07 V_hig
+ 2.770010000e-07 V_hig
+ 2.771000000e-07 V_hig
+ 2.771010000e-07 V_hig
+ 2.772000000e-07 V_hig
+ 2.772010000e-07 V_hig
+ 2.773000000e-07 V_hig
+ 2.773010000e-07 V_hig
+ 2.774000000e-07 V_hig
+ 2.774010000e-07 V_hig
+ 2.775000000e-07 V_hig
+ 2.775010000e-07 V_hig
+ 2.776000000e-07 V_hig
+ 2.776010000e-07 V_hig
+ 2.777000000e-07 V_hig
+ 2.777010000e-07 V_hig
+ 2.778000000e-07 V_hig
+ 2.778010000e-07 V_hig
+ 2.779000000e-07 V_hig
+ 2.779010000e-07 V_hig
+ 2.780000000e-07 V_hig
+ 2.780010000e-07 V_hig
+ 2.781000000e-07 V_hig
+ 2.781010000e-07 V_hig
+ 2.782000000e-07 V_hig
+ 2.782010000e-07 V_hig
+ 2.783000000e-07 V_hig
+ 2.783010000e-07 V_hig
+ 2.784000000e-07 V_hig
+ 2.784010000e-07 V_hig
+ 2.785000000e-07 V_hig
+ 2.785010000e-07 V_hig
+ 2.786000000e-07 V_hig
+ 2.786010000e-07 V_hig
+ 2.787000000e-07 V_hig
+ 2.787010000e-07 V_hig
+ 2.788000000e-07 V_hig
+ 2.788010000e-07 V_hig
+ 2.789000000e-07 V_hig
+ 2.789010000e-07 V_low
+ 2.790000000e-07 V_low
+ 2.790010000e-07 V_low
+ 2.791000000e-07 V_low
+ 2.791010000e-07 V_low
+ 2.792000000e-07 V_low
+ 2.792010000e-07 V_low
+ 2.793000000e-07 V_low
+ 2.793010000e-07 V_low
+ 2.794000000e-07 V_low
+ 2.794010000e-07 V_low
+ 2.795000000e-07 V_low
+ 2.795010000e-07 V_low
+ 2.796000000e-07 V_low
+ 2.796010000e-07 V_low
+ 2.797000000e-07 V_low
+ 2.797010000e-07 V_low
+ 2.798000000e-07 V_low
+ 2.798010000e-07 V_low
+ 2.799000000e-07 V_low
+ 2.799010000e-07 V_hig
+ 2.800000000e-07 V_hig
+ 2.800010000e-07 V_hig
+ 2.801000000e-07 V_hig
+ 2.801010000e-07 V_hig
+ 2.802000000e-07 V_hig
+ 2.802010000e-07 V_hig
+ 2.803000000e-07 V_hig
+ 2.803010000e-07 V_hig
+ 2.804000000e-07 V_hig
+ 2.804010000e-07 V_hig
+ 2.805000000e-07 V_hig
+ 2.805010000e-07 V_hig
+ 2.806000000e-07 V_hig
+ 2.806010000e-07 V_hig
+ 2.807000000e-07 V_hig
+ 2.807010000e-07 V_hig
+ 2.808000000e-07 V_hig
+ 2.808010000e-07 V_hig
+ 2.809000000e-07 V_hig
+ 2.809010000e-07 V_low
+ 2.810000000e-07 V_low
+ 2.810010000e-07 V_low
+ 2.811000000e-07 V_low
+ 2.811010000e-07 V_low
+ 2.812000000e-07 V_low
+ 2.812010000e-07 V_low
+ 2.813000000e-07 V_low
+ 2.813010000e-07 V_low
+ 2.814000000e-07 V_low
+ 2.814010000e-07 V_low
+ 2.815000000e-07 V_low
+ 2.815010000e-07 V_low
+ 2.816000000e-07 V_low
+ 2.816010000e-07 V_low
+ 2.817000000e-07 V_low
+ 2.817010000e-07 V_low
+ 2.818000000e-07 V_low
+ 2.818010000e-07 V_low
+ 2.819000000e-07 V_low
+ 2.819010000e-07 V_low
+ 2.820000000e-07 V_low
+ 2.820010000e-07 V_low
+ 2.821000000e-07 V_low
+ 2.821010000e-07 V_low
+ 2.822000000e-07 V_low
+ 2.822010000e-07 V_low
+ 2.823000000e-07 V_low
+ 2.823010000e-07 V_low
+ 2.824000000e-07 V_low
+ 2.824010000e-07 V_low
+ 2.825000000e-07 V_low
+ 2.825010000e-07 V_low
+ 2.826000000e-07 V_low
+ 2.826010000e-07 V_low
+ 2.827000000e-07 V_low
+ 2.827010000e-07 V_low
+ 2.828000000e-07 V_low
+ 2.828010000e-07 V_low
+ 2.829000000e-07 V_low
+ 2.829010000e-07 V_hig
+ 2.830000000e-07 V_hig
+ 2.830010000e-07 V_hig
+ 2.831000000e-07 V_hig
+ 2.831010000e-07 V_hig
+ 2.832000000e-07 V_hig
+ 2.832010000e-07 V_hig
+ 2.833000000e-07 V_hig
+ 2.833010000e-07 V_hig
+ 2.834000000e-07 V_hig
+ 2.834010000e-07 V_hig
+ 2.835000000e-07 V_hig
+ 2.835010000e-07 V_hig
+ 2.836000000e-07 V_hig
+ 2.836010000e-07 V_hig
+ 2.837000000e-07 V_hig
+ 2.837010000e-07 V_hig
+ 2.838000000e-07 V_hig
+ 2.838010000e-07 V_hig
+ 2.839000000e-07 V_hig
+ 2.839010000e-07 V_low
+ 2.840000000e-07 V_low
+ 2.840010000e-07 V_low
+ 2.841000000e-07 V_low
+ 2.841010000e-07 V_low
+ 2.842000000e-07 V_low
+ 2.842010000e-07 V_low
+ 2.843000000e-07 V_low
+ 2.843010000e-07 V_low
+ 2.844000000e-07 V_low
+ 2.844010000e-07 V_low
+ 2.845000000e-07 V_low
+ 2.845010000e-07 V_low
+ 2.846000000e-07 V_low
+ 2.846010000e-07 V_low
+ 2.847000000e-07 V_low
+ 2.847010000e-07 V_low
+ 2.848000000e-07 V_low
+ 2.848010000e-07 V_low
+ 2.849000000e-07 V_low
+ 2.849010000e-07 V_low
+ 2.850000000e-07 V_low
+ 2.850010000e-07 V_low
+ 2.851000000e-07 V_low
+ 2.851010000e-07 V_low
+ 2.852000000e-07 V_low
+ 2.852010000e-07 V_low
+ 2.853000000e-07 V_low
+ 2.853010000e-07 V_low
+ 2.854000000e-07 V_low
+ 2.854010000e-07 V_low
+ 2.855000000e-07 V_low
+ 2.855010000e-07 V_low
+ 2.856000000e-07 V_low
+ 2.856010000e-07 V_low
+ 2.857000000e-07 V_low
+ 2.857010000e-07 V_low
+ 2.858000000e-07 V_low
+ 2.858010000e-07 V_low
+ 2.859000000e-07 V_low
+ 2.859010000e-07 V_hig
+ 2.860000000e-07 V_hig
+ 2.860010000e-07 V_hig
+ 2.861000000e-07 V_hig
+ 2.861010000e-07 V_hig
+ 2.862000000e-07 V_hig
+ 2.862010000e-07 V_hig
+ 2.863000000e-07 V_hig
+ 2.863010000e-07 V_hig
+ 2.864000000e-07 V_hig
+ 2.864010000e-07 V_hig
+ 2.865000000e-07 V_hig
+ 2.865010000e-07 V_hig
+ 2.866000000e-07 V_hig
+ 2.866010000e-07 V_hig
+ 2.867000000e-07 V_hig
+ 2.867010000e-07 V_hig
+ 2.868000000e-07 V_hig
+ 2.868010000e-07 V_hig
+ 2.869000000e-07 V_hig
+ 2.869010000e-07 V_hig
+ 2.870000000e-07 V_hig
+ 2.870010000e-07 V_hig
+ 2.871000000e-07 V_hig
+ 2.871010000e-07 V_hig
+ 2.872000000e-07 V_hig
+ 2.872010000e-07 V_hig
+ 2.873000000e-07 V_hig
+ 2.873010000e-07 V_hig
+ 2.874000000e-07 V_hig
+ 2.874010000e-07 V_hig
+ 2.875000000e-07 V_hig
+ 2.875010000e-07 V_hig
+ 2.876000000e-07 V_hig
+ 2.876010000e-07 V_hig
+ 2.877000000e-07 V_hig
+ 2.877010000e-07 V_hig
+ 2.878000000e-07 V_hig
+ 2.878010000e-07 V_hig
+ 2.879000000e-07 V_hig
+ 2.879010000e-07 V_hig
+ 2.880000000e-07 V_hig
+ 2.880010000e-07 V_hig
+ 2.881000000e-07 V_hig
+ 2.881010000e-07 V_hig
+ 2.882000000e-07 V_hig
+ 2.882010000e-07 V_hig
+ 2.883000000e-07 V_hig
+ 2.883010000e-07 V_hig
+ 2.884000000e-07 V_hig
+ 2.884010000e-07 V_hig
+ 2.885000000e-07 V_hig
+ 2.885010000e-07 V_hig
+ 2.886000000e-07 V_hig
+ 2.886010000e-07 V_hig
+ 2.887000000e-07 V_hig
+ 2.887010000e-07 V_hig
+ 2.888000000e-07 V_hig
+ 2.888010000e-07 V_hig
+ 2.889000000e-07 V_hig
+ 2.889010000e-07 V_hig
+ 2.890000000e-07 V_hig
+ 2.890010000e-07 V_hig
+ 2.891000000e-07 V_hig
+ 2.891010000e-07 V_hig
+ 2.892000000e-07 V_hig
+ 2.892010000e-07 V_hig
+ 2.893000000e-07 V_hig
+ 2.893010000e-07 V_hig
+ 2.894000000e-07 V_hig
+ 2.894010000e-07 V_hig
+ 2.895000000e-07 V_hig
+ 2.895010000e-07 V_hig
+ 2.896000000e-07 V_hig
+ 2.896010000e-07 V_hig
+ 2.897000000e-07 V_hig
+ 2.897010000e-07 V_hig
+ 2.898000000e-07 V_hig
+ 2.898010000e-07 V_hig
+ 2.899000000e-07 V_hig
+ 2.899010000e-07 V_hig
+ 2.900000000e-07 V_hig
+ 2.900010000e-07 V_hig
+ 2.901000000e-07 V_hig
+ 2.901010000e-07 V_hig
+ 2.902000000e-07 V_hig
+ 2.902010000e-07 V_hig
+ 2.903000000e-07 V_hig
+ 2.903010000e-07 V_hig
+ 2.904000000e-07 V_hig
+ 2.904010000e-07 V_hig
+ 2.905000000e-07 V_hig
+ 2.905010000e-07 V_hig
+ 2.906000000e-07 V_hig
+ 2.906010000e-07 V_hig
+ 2.907000000e-07 V_hig
+ 2.907010000e-07 V_hig
+ 2.908000000e-07 V_hig
+ 2.908010000e-07 V_hig
+ 2.909000000e-07 V_hig
+ 2.909010000e-07 V_low
+ 2.910000000e-07 V_low
+ 2.910010000e-07 V_low
+ 2.911000000e-07 V_low
+ 2.911010000e-07 V_low
+ 2.912000000e-07 V_low
+ 2.912010000e-07 V_low
+ 2.913000000e-07 V_low
+ 2.913010000e-07 V_low
+ 2.914000000e-07 V_low
+ 2.914010000e-07 V_low
+ 2.915000000e-07 V_low
+ 2.915010000e-07 V_low
+ 2.916000000e-07 V_low
+ 2.916010000e-07 V_low
+ 2.917000000e-07 V_low
+ 2.917010000e-07 V_low
+ 2.918000000e-07 V_low
+ 2.918010000e-07 V_low
+ 2.919000000e-07 V_low
+ 2.919010000e-07 V_low
+ 2.920000000e-07 V_low
+ 2.920010000e-07 V_low
+ 2.921000000e-07 V_low
+ 2.921010000e-07 V_low
+ 2.922000000e-07 V_low
+ 2.922010000e-07 V_low
+ 2.923000000e-07 V_low
+ 2.923010000e-07 V_low
+ 2.924000000e-07 V_low
+ 2.924010000e-07 V_low
+ 2.925000000e-07 V_low
+ 2.925010000e-07 V_low
+ 2.926000000e-07 V_low
+ 2.926010000e-07 V_low
+ 2.927000000e-07 V_low
+ 2.927010000e-07 V_low
+ 2.928000000e-07 V_low
+ 2.928010000e-07 V_low
+ 2.929000000e-07 V_low
+ 2.929010000e-07 V_hig
+ 2.930000000e-07 V_hig
+ 2.930010000e-07 V_hig
+ 2.931000000e-07 V_hig
+ 2.931010000e-07 V_hig
+ 2.932000000e-07 V_hig
+ 2.932010000e-07 V_hig
+ 2.933000000e-07 V_hig
+ 2.933010000e-07 V_hig
+ 2.934000000e-07 V_hig
+ 2.934010000e-07 V_hig
+ 2.935000000e-07 V_hig
+ 2.935010000e-07 V_hig
+ 2.936000000e-07 V_hig
+ 2.936010000e-07 V_hig
+ 2.937000000e-07 V_hig
+ 2.937010000e-07 V_hig
+ 2.938000000e-07 V_hig
+ 2.938010000e-07 V_hig
+ 2.939000000e-07 V_hig
+ 2.939010000e-07 V_low
+ 2.940000000e-07 V_low
+ 2.940010000e-07 V_low
+ 2.941000000e-07 V_low
+ 2.941010000e-07 V_low
+ 2.942000000e-07 V_low
+ 2.942010000e-07 V_low
+ 2.943000000e-07 V_low
+ 2.943010000e-07 V_low
+ 2.944000000e-07 V_low
+ 2.944010000e-07 V_low
+ 2.945000000e-07 V_low
+ 2.945010000e-07 V_low
+ 2.946000000e-07 V_low
+ 2.946010000e-07 V_low
+ 2.947000000e-07 V_low
+ 2.947010000e-07 V_low
+ 2.948000000e-07 V_low
+ 2.948010000e-07 V_low
+ 2.949000000e-07 V_low
+ 2.949010000e-07 V_low
+ 2.950000000e-07 V_low
+ 2.950010000e-07 V_low
+ 2.951000000e-07 V_low
+ 2.951010000e-07 V_low
+ 2.952000000e-07 V_low
+ 2.952010000e-07 V_low
+ 2.953000000e-07 V_low
+ 2.953010000e-07 V_low
+ 2.954000000e-07 V_low
+ 2.954010000e-07 V_low
+ 2.955000000e-07 V_low
+ 2.955010000e-07 V_low
+ 2.956000000e-07 V_low
+ 2.956010000e-07 V_low
+ 2.957000000e-07 V_low
+ 2.957010000e-07 V_low
+ 2.958000000e-07 V_low
+ 2.958010000e-07 V_low
+ 2.959000000e-07 V_low
+ 2.959010000e-07 V_hig
+ 2.960000000e-07 V_hig
+ 2.960010000e-07 V_hig
+ 2.961000000e-07 V_hig
+ 2.961010000e-07 V_hig
+ 2.962000000e-07 V_hig
+ 2.962010000e-07 V_hig
+ 2.963000000e-07 V_hig
+ 2.963010000e-07 V_hig
+ 2.964000000e-07 V_hig
+ 2.964010000e-07 V_hig
+ 2.965000000e-07 V_hig
+ 2.965010000e-07 V_hig
+ 2.966000000e-07 V_hig
+ 2.966010000e-07 V_hig
+ 2.967000000e-07 V_hig
+ 2.967010000e-07 V_hig
+ 2.968000000e-07 V_hig
+ 2.968010000e-07 V_hig
+ 2.969000000e-07 V_hig
+ 2.969010000e-07 V_hig
+ 2.970000000e-07 V_hig
+ 2.970010000e-07 V_hig
+ 2.971000000e-07 V_hig
+ 2.971010000e-07 V_hig
+ 2.972000000e-07 V_hig
+ 2.972010000e-07 V_hig
+ 2.973000000e-07 V_hig
+ 2.973010000e-07 V_hig
+ 2.974000000e-07 V_hig
+ 2.974010000e-07 V_hig
+ 2.975000000e-07 V_hig
+ 2.975010000e-07 V_hig
+ 2.976000000e-07 V_hig
+ 2.976010000e-07 V_hig
+ 2.977000000e-07 V_hig
+ 2.977010000e-07 V_hig
+ 2.978000000e-07 V_hig
+ 2.978010000e-07 V_hig
+ 2.979000000e-07 V_hig
+ 2.979010000e-07 V_low
+ 2.980000000e-07 V_low
+ 2.980010000e-07 V_low
+ 2.981000000e-07 V_low
+ 2.981010000e-07 V_low
+ 2.982000000e-07 V_low
+ 2.982010000e-07 V_low
+ 2.983000000e-07 V_low
+ 2.983010000e-07 V_low
+ 2.984000000e-07 V_low
+ 2.984010000e-07 V_low
+ 2.985000000e-07 V_low
+ 2.985010000e-07 V_low
+ 2.986000000e-07 V_low
+ 2.986010000e-07 V_low
+ 2.987000000e-07 V_low
+ 2.987010000e-07 V_low
+ 2.988000000e-07 V_low
+ 2.988010000e-07 V_low
+ 2.989000000e-07 V_low
+ 2.989010000e-07 V_hig
+ 2.990000000e-07 V_hig
+ 2.990010000e-07 V_hig
+ 2.991000000e-07 V_hig
+ 2.991010000e-07 V_hig
+ 2.992000000e-07 V_hig
+ 2.992010000e-07 V_hig
+ 2.993000000e-07 V_hig
+ 2.993010000e-07 V_hig
+ 2.994000000e-07 V_hig
+ 2.994010000e-07 V_hig
+ 2.995000000e-07 V_hig
+ 2.995010000e-07 V_hig
+ 2.996000000e-07 V_hig
+ 2.996010000e-07 V_hig
+ 2.997000000e-07 V_hig
+ 2.997010000e-07 V_hig
+ 2.998000000e-07 V_hig
+ 2.998010000e-07 V_hig
+ 2.999000000e-07 V_hig
+ 2.999010000e-07 V_hig
+ 3.000000000e-07 V_hig
+ 3.000010000e-07 V_hig
+ 3.001000000e-07 V_hig
+ 3.001010000e-07 V_hig
+ 3.002000000e-07 V_hig
+ 3.002010000e-07 V_hig
+ 3.003000000e-07 V_hig
+ 3.003010000e-07 V_hig
+ 3.004000000e-07 V_hig
+ 3.004010000e-07 V_hig
+ 3.005000000e-07 V_hig
+ 3.005010000e-07 V_hig
+ 3.006000000e-07 V_hig
+ 3.006010000e-07 V_hig
+ 3.007000000e-07 V_hig
+ 3.007010000e-07 V_hig
+ 3.008000000e-07 V_hig
+ 3.008010000e-07 V_hig
+ 3.009000000e-07 V_hig
+ 3.009010000e-07 V_low
+ 3.010000000e-07 V_low
+ 3.010010000e-07 V_low
+ 3.011000000e-07 V_low
+ 3.011010000e-07 V_low
+ 3.012000000e-07 V_low
+ 3.012010000e-07 V_low
+ 3.013000000e-07 V_low
+ 3.013010000e-07 V_low
+ 3.014000000e-07 V_low
+ 3.014010000e-07 V_low
+ 3.015000000e-07 V_low
+ 3.015010000e-07 V_low
+ 3.016000000e-07 V_low
+ 3.016010000e-07 V_low
+ 3.017000000e-07 V_low
+ 3.017010000e-07 V_low
+ 3.018000000e-07 V_low
+ 3.018010000e-07 V_low
+ 3.019000000e-07 V_low
+ 3.019010000e-07 V_hig
+ 3.020000000e-07 V_hig
+ 3.020010000e-07 V_hig
+ 3.021000000e-07 V_hig
+ 3.021010000e-07 V_hig
+ 3.022000000e-07 V_hig
+ 3.022010000e-07 V_hig
+ 3.023000000e-07 V_hig
+ 3.023010000e-07 V_hig
+ 3.024000000e-07 V_hig
+ 3.024010000e-07 V_hig
+ 3.025000000e-07 V_hig
+ 3.025010000e-07 V_hig
+ 3.026000000e-07 V_hig
+ 3.026010000e-07 V_hig
+ 3.027000000e-07 V_hig
+ 3.027010000e-07 V_hig
+ 3.028000000e-07 V_hig
+ 3.028010000e-07 V_hig
+ 3.029000000e-07 V_hig
+ 3.029010000e-07 V_low
+ 3.030000000e-07 V_low
+ 3.030010000e-07 V_low
+ 3.031000000e-07 V_low
+ 3.031010000e-07 V_low
+ 3.032000000e-07 V_low
+ 3.032010000e-07 V_low
+ 3.033000000e-07 V_low
+ 3.033010000e-07 V_low
+ 3.034000000e-07 V_low
+ 3.034010000e-07 V_low
+ 3.035000000e-07 V_low
+ 3.035010000e-07 V_low
+ 3.036000000e-07 V_low
+ 3.036010000e-07 V_low
+ 3.037000000e-07 V_low
+ 3.037010000e-07 V_low
+ 3.038000000e-07 V_low
+ 3.038010000e-07 V_low
+ 3.039000000e-07 V_low
+ 3.039010000e-07 V_low
+ 3.040000000e-07 V_low
+ 3.040010000e-07 V_low
+ 3.041000000e-07 V_low
+ 3.041010000e-07 V_low
+ 3.042000000e-07 V_low
+ 3.042010000e-07 V_low
+ 3.043000000e-07 V_low
+ 3.043010000e-07 V_low
+ 3.044000000e-07 V_low
+ 3.044010000e-07 V_low
+ 3.045000000e-07 V_low
+ 3.045010000e-07 V_low
+ 3.046000000e-07 V_low
+ 3.046010000e-07 V_low
+ 3.047000000e-07 V_low
+ 3.047010000e-07 V_low
+ 3.048000000e-07 V_low
+ 3.048010000e-07 V_low
+ 3.049000000e-07 V_low
+ 3.049010000e-07 V_low
+ 3.050000000e-07 V_low
+ 3.050010000e-07 V_low
+ 3.051000000e-07 V_low
+ 3.051010000e-07 V_low
+ 3.052000000e-07 V_low
+ 3.052010000e-07 V_low
+ 3.053000000e-07 V_low
+ 3.053010000e-07 V_low
+ 3.054000000e-07 V_low
+ 3.054010000e-07 V_low
+ 3.055000000e-07 V_low
+ 3.055010000e-07 V_low
+ 3.056000000e-07 V_low
+ 3.056010000e-07 V_low
+ 3.057000000e-07 V_low
+ 3.057010000e-07 V_low
+ 3.058000000e-07 V_low
+ 3.058010000e-07 V_low
+ 3.059000000e-07 V_low
+ 3.059010000e-07 V_hig
+ 3.060000000e-07 V_hig
+ 3.060010000e-07 V_hig
+ 3.061000000e-07 V_hig
+ 3.061010000e-07 V_hig
+ 3.062000000e-07 V_hig
+ 3.062010000e-07 V_hig
+ 3.063000000e-07 V_hig
+ 3.063010000e-07 V_hig
+ 3.064000000e-07 V_hig
+ 3.064010000e-07 V_hig
+ 3.065000000e-07 V_hig
+ 3.065010000e-07 V_hig
+ 3.066000000e-07 V_hig
+ 3.066010000e-07 V_hig
+ 3.067000000e-07 V_hig
+ 3.067010000e-07 V_hig
+ 3.068000000e-07 V_hig
+ 3.068010000e-07 V_hig
+ 3.069000000e-07 V_hig
+ 3.069010000e-07 V_hig
+ 3.070000000e-07 V_hig
+ 3.070010000e-07 V_hig
+ 3.071000000e-07 V_hig
+ 3.071010000e-07 V_hig
+ 3.072000000e-07 V_hig
+ 3.072010000e-07 V_hig
+ 3.073000000e-07 V_hig
+ 3.073010000e-07 V_hig
+ 3.074000000e-07 V_hig
+ 3.074010000e-07 V_hig
+ 3.075000000e-07 V_hig
+ 3.075010000e-07 V_hig
+ 3.076000000e-07 V_hig
+ 3.076010000e-07 V_hig
+ 3.077000000e-07 V_hig
+ 3.077010000e-07 V_hig
+ 3.078000000e-07 V_hig
+ 3.078010000e-07 V_hig
+ 3.079000000e-07 V_hig
+ 3.079010000e-07 V_low
+ 3.080000000e-07 V_low
+ 3.080010000e-07 V_low
+ 3.081000000e-07 V_low
+ 3.081010000e-07 V_low
+ 3.082000000e-07 V_low
+ 3.082010000e-07 V_low
+ 3.083000000e-07 V_low
+ 3.083010000e-07 V_low
+ 3.084000000e-07 V_low
+ 3.084010000e-07 V_low
+ 3.085000000e-07 V_low
+ 3.085010000e-07 V_low
+ 3.086000000e-07 V_low
+ 3.086010000e-07 V_low
+ 3.087000000e-07 V_low
+ 3.087010000e-07 V_low
+ 3.088000000e-07 V_low
+ 3.088010000e-07 V_low
+ 3.089000000e-07 V_low
+ 3.089010000e-07 V_low
+ 3.090000000e-07 V_low
+ 3.090010000e-07 V_low
+ 3.091000000e-07 V_low
+ 3.091010000e-07 V_low
+ 3.092000000e-07 V_low
+ 3.092010000e-07 V_low
+ 3.093000000e-07 V_low
+ 3.093010000e-07 V_low
+ 3.094000000e-07 V_low
+ 3.094010000e-07 V_low
+ 3.095000000e-07 V_low
+ 3.095010000e-07 V_low
+ 3.096000000e-07 V_low
+ 3.096010000e-07 V_low
+ 3.097000000e-07 V_low
+ 3.097010000e-07 V_low
+ 3.098000000e-07 V_low
+ 3.098010000e-07 V_low
+ 3.099000000e-07 V_low
+ 3.099010000e-07 V_low
+ 3.100000000e-07 V_low
+ 3.100010000e-07 V_low
+ 3.101000000e-07 V_low
+ 3.101010000e-07 V_low
+ 3.102000000e-07 V_low
+ 3.102010000e-07 V_low
+ 3.103000000e-07 V_low
+ 3.103010000e-07 V_low
+ 3.104000000e-07 V_low
+ 3.104010000e-07 V_low
+ 3.105000000e-07 V_low
+ 3.105010000e-07 V_low
+ 3.106000000e-07 V_low
+ 3.106010000e-07 V_low
+ 3.107000000e-07 V_low
+ 3.107010000e-07 V_low
+ 3.108000000e-07 V_low
+ 3.108010000e-07 V_low
+ 3.109000000e-07 V_low
+ 3.109010000e-07 V_low
+ 3.110000000e-07 V_low
+ 3.110010000e-07 V_low
+ 3.111000000e-07 V_low
+ 3.111010000e-07 V_low
+ 3.112000000e-07 V_low
+ 3.112010000e-07 V_low
+ 3.113000000e-07 V_low
+ 3.113010000e-07 V_low
+ 3.114000000e-07 V_low
+ 3.114010000e-07 V_low
+ 3.115000000e-07 V_low
+ 3.115010000e-07 V_low
+ 3.116000000e-07 V_low
+ 3.116010000e-07 V_low
+ 3.117000000e-07 V_low
+ 3.117010000e-07 V_low
+ 3.118000000e-07 V_low
+ 3.118010000e-07 V_low
+ 3.119000000e-07 V_low
+ 3.119010000e-07 V_low
+ 3.120000000e-07 V_low
+ 3.120010000e-07 V_low
+ 3.121000000e-07 V_low
+ 3.121010000e-07 V_low
+ 3.122000000e-07 V_low
+ 3.122010000e-07 V_low
+ 3.123000000e-07 V_low
+ 3.123010000e-07 V_low
+ 3.124000000e-07 V_low
+ 3.124010000e-07 V_low
+ 3.125000000e-07 V_low
+ 3.125010000e-07 V_low
+ 3.126000000e-07 V_low
+ 3.126010000e-07 V_low
+ 3.127000000e-07 V_low
+ 3.127010000e-07 V_low
+ 3.128000000e-07 V_low
+ 3.128010000e-07 V_low
+ 3.129000000e-07 V_low
+ 3.129010000e-07 V_low
+ 3.130000000e-07 V_low
+ 3.130010000e-07 V_low
+ 3.131000000e-07 V_low
+ 3.131010000e-07 V_low
+ 3.132000000e-07 V_low
+ 3.132010000e-07 V_low
+ 3.133000000e-07 V_low
+ 3.133010000e-07 V_low
+ 3.134000000e-07 V_low
+ 3.134010000e-07 V_low
+ 3.135000000e-07 V_low
+ 3.135010000e-07 V_low
+ 3.136000000e-07 V_low
+ 3.136010000e-07 V_low
+ 3.137000000e-07 V_low
+ 3.137010000e-07 V_low
+ 3.138000000e-07 V_low
+ 3.138010000e-07 V_low
+ 3.139000000e-07 V_low
+ 3.139010000e-07 V_low
+ 3.140000000e-07 V_low
+ 3.140010000e-07 V_low
+ 3.141000000e-07 V_low
+ 3.141010000e-07 V_low
+ 3.142000000e-07 V_low
+ 3.142010000e-07 V_low
+ 3.143000000e-07 V_low
+ 3.143010000e-07 V_low
+ 3.144000000e-07 V_low
+ 3.144010000e-07 V_low
+ 3.145000000e-07 V_low
+ 3.145010000e-07 V_low
+ 3.146000000e-07 V_low
+ 3.146010000e-07 V_low
+ 3.147000000e-07 V_low
+ 3.147010000e-07 V_low
+ 3.148000000e-07 V_low
+ 3.148010000e-07 V_low
+ 3.149000000e-07 V_low
+ 3.149010000e-07 V_low
+ 3.150000000e-07 V_low
+ 3.150010000e-07 V_low
+ 3.151000000e-07 V_low
+ 3.151010000e-07 V_low
+ 3.152000000e-07 V_low
+ 3.152010000e-07 V_low
+ 3.153000000e-07 V_low
+ 3.153010000e-07 V_low
+ 3.154000000e-07 V_low
+ 3.154010000e-07 V_low
+ 3.155000000e-07 V_low
+ 3.155010000e-07 V_low
+ 3.156000000e-07 V_low
+ 3.156010000e-07 V_low
+ 3.157000000e-07 V_low
+ 3.157010000e-07 V_low
+ 3.158000000e-07 V_low
+ 3.158010000e-07 V_low
+ 3.159000000e-07 V_low
+ 3.159010000e-07 V_hig
+ 3.160000000e-07 V_hig
+ 3.160010000e-07 V_hig
+ 3.161000000e-07 V_hig
+ 3.161010000e-07 V_hig
+ 3.162000000e-07 V_hig
+ 3.162010000e-07 V_hig
+ 3.163000000e-07 V_hig
+ 3.163010000e-07 V_hig
+ 3.164000000e-07 V_hig
+ 3.164010000e-07 V_hig
+ 3.165000000e-07 V_hig
+ 3.165010000e-07 V_hig
+ 3.166000000e-07 V_hig
+ 3.166010000e-07 V_hig
+ 3.167000000e-07 V_hig
+ 3.167010000e-07 V_hig
+ 3.168000000e-07 V_hig
+ 3.168010000e-07 V_hig
+ 3.169000000e-07 V_hig
+ 3.169010000e-07 V_low
+ 3.170000000e-07 V_low
+ 3.170010000e-07 V_low
+ 3.171000000e-07 V_low
+ 3.171010000e-07 V_low
+ 3.172000000e-07 V_low
+ 3.172010000e-07 V_low
+ 3.173000000e-07 V_low
+ 3.173010000e-07 V_low
+ 3.174000000e-07 V_low
+ 3.174010000e-07 V_low
+ 3.175000000e-07 V_low
+ 3.175010000e-07 V_low
+ 3.176000000e-07 V_low
+ 3.176010000e-07 V_low
+ 3.177000000e-07 V_low
+ 3.177010000e-07 V_low
+ 3.178000000e-07 V_low
+ 3.178010000e-07 V_low
+ 3.179000000e-07 V_low
+ 3.179010000e-07 V_hig
+ 3.180000000e-07 V_hig
+ 3.180010000e-07 V_hig
+ 3.181000000e-07 V_hig
+ 3.181010000e-07 V_hig
+ 3.182000000e-07 V_hig
+ 3.182010000e-07 V_hig
+ 3.183000000e-07 V_hig
+ 3.183010000e-07 V_hig
+ 3.184000000e-07 V_hig
+ 3.184010000e-07 V_hig
+ 3.185000000e-07 V_hig
+ 3.185010000e-07 V_hig
+ 3.186000000e-07 V_hig
+ 3.186010000e-07 V_hig
+ 3.187000000e-07 V_hig
+ 3.187010000e-07 V_hig
+ 3.188000000e-07 V_hig
+ 3.188010000e-07 V_hig
+ 3.189000000e-07 V_hig
+ 3.189010000e-07 V_low
+ 3.190000000e-07 V_low
+ 3.190010000e-07 V_low
+ 3.191000000e-07 V_low
+ 3.191010000e-07 V_low
+ 3.192000000e-07 V_low
+ 3.192010000e-07 V_low
+ 3.193000000e-07 V_low
+ 3.193010000e-07 V_low
+ 3.194000000e-07 V_low
+ 3.194010000e-07 V_low
+ 3.195000000e-07 V_low
+ 3.195010000e-07 V_low
+ 3.196000000e-07 V_low
+ 3.196010000e-07 V_low
+ 3.197000000e-07 V_low
+ 3.197010000e-07 V_low
+ 3.198000000e-07 V_low
+ 3.198010000e-07 V_low
+ 3.199000000e-07 V_low
+ 3.199010000e-07 V_hig
+ 3.200000000e-07 V_hig
+ 3.200010000e-07 V_hig
+ 3.201000000e-07 V_hig
+ 3.201010000e-07 V_hig
+ 3.202000000e-07 V_hig
+ 3.202010000e-07 V_hig
+ 3.203000000e-07 V_hig
+ 3.203010000e-07 V_hig
+ 3.204000000e-07 V_hig
+ 3.204010000e-07 V_hig
+ 3.205000000e-07 V_hig
+ 3.205010000e-07 V_hig
+ 3.206000000e-07 V_hig
+ 3.206010000e-07 V_hig
+ 3.207000000e-07 V_hig
+ 3.207010000e-07 V_hig
+ 3.208000000e-07 V_hig
+ 3.208010000e-07 V_hig
+ 3.209000000e-07 V_hig
+ 3.209010000e-07 V_hig
+ 3.210000000e-07 V_hig
+ 3.210010000e-07 V_hig
+ 3.211000000e-07 V_hig
+ 3.211010000e-07 V_hig
+ 3.212000000e-07 V_hig
+ 3.212010000e-07 V_hig
+ 3.213000000e-07 V_hig
+ 3.213010000e-07 V_hig
+ 3.214000000e-07 V_hig
+ 3.214010000e-07 V_hig
+ 3.215000000e-07 V_hig
+ 3.215010000e-07 V_hig
+ 3.216000000e-07 V_hig
+ 3.216010000e-07 V_hig
+ 3.217000000e-07 V_hig
+ 3.217010000e-07 V_hig
+ 3.218000000e-07 V_hig
+ 3.218010000e-07 V_hig
+ 3.219000000e-07 V_hig
+ 3.219010000e-07 V_hig
+ 3.220000000e-07 V_hig
+ 3.220010000e-07 V_hig
+ 3.221000000e-07 V_hig
+ 3.221010000e-07 V_hig
+ 3.222000000e-07 V_hig
+ 3.222010000e-07 V_hig
+ 3.223000000e-07 V_hig
+ 3.223010000e-07 V_hig
+ 3.224000000e-07 V_hig
+ 3.224010000e-07 V_hig
+ 3.225000000e-07 V_hig
+ 3.225010000e-07 V_hig
+ 3.226000000e-07 V_hig
+ 3.226010000e-07 V_hig
+ 3.227000000e-07 V_hig
+ 3.227010000e-07 V_hig
+ 3.228000000e-07 V_hig
+ 3.228010000e-07 V_hig
+ 3.229000000e-07 V_hig
+ 3.229010000e-07 V_low
+ 3.230000000e-07 V_low
+ 3.230010000e-07 V_low
+ 3.231000000e-07 V_low
+ 3.231010000e-07 V_low
+ 3.232000000e-07 V_low
+ 3.232010000e-07 V_low
+ 3.233000000e-07 V_low
+ 3.233010000e-07 V_low
+ 3.234000000e-07 V_low
+ 3.234010000e-07 V_low
+ 3.235000000e-07 V_low
+ 3.235010000e-07 V_low
+ 3.236000000e-07 V_low
+ 3.236010000e-07 V_low
+ 3.237000000e-07 V_low
+ 3.237010000e-07 V_low
+ 3.238000000e-07 V_low
+ 3.238010000e-07 V_low
+ 3.239000000e-07 V_low
+ 3.239010000e-07 V_hig
+ 3.240000000e-07 V_hig
+ 3.240010000e-07 V_hig
+ 3.241000000e-07 V_hig
+ 3.241010000e-07 V_hig
+ 3.242000000e-07 V_hig
+ 3.242010000e-07 V_hig
+ 3.243000000e-07 V_hig
+ 3.243010000e-07 V_hig
+ 3.244000000e-07 V_hig
+ 3.244010000e-07 V_hig
+ 3.245000000e-07 V_hig
+ 3.245010000e-07 V_hig
+ 3.246000000e-07 V_hig
+ 3.246010000e-07 V_hig
+ 3.247000000e-07 V_hig
+ 3.247010000e-07 V_hig
+ 3.248000000e-07 V_hig
+ 3.248010000e-07 V_hig
+ 3.249000000e-07 V_hig
+ 3.249010000e-07 V_hig
+ 3.250000000e-07 V_hig
+ 3.250010000e-07 V_hig
+ 3.251000000e-07 V_hig
+ 3.251010000e-07 V_hig
+ 3.252000000e-07 V_hig
+ 3.252010000e-07 V_hig
+ 3.253000000e-07 V_hig
+ 3.253010000e-07 V_hig
+ 3.254000000e-07 V_hig
+ 3.254010000e-07 V_hig
+ 3.255000000e-07 V_hig
+ 3.255010000e-07 V_hig
+ 3.256000000e-07 V_hig
+ 3.256010000e-07 V_hig
+ 3.257000000e-07 V_hig
+ 3.257010000e-07 V_hig
+ 3.258000000e-07 V_hig
+ 3.258010000e-07 V_hig
+ 3.259000000e-07 V_hig
+ 3.259010000e-07 V_low
+ 3.260000000e-07 V_low
+ 3.260010000e-07 V_low
+ 3.261000000e-07 V_low
+ 3.261010000e-07 V_low
+ 3.262000000e-07 V_low
+ 3.262010000e-07 V_low
+ 3.263000000e-07 V_low
+ 3.263010000e-07 V_low
+ 3.264000000e-07 V_low
+ 3.264010000e-07 V_low
+ 3.265000000e-07 V_low
+ 3.265010000e-07 V_low
+ 3.266000000e-07 V_low
+ 3.266010000e-07 V_low
+ 3.267000000e-07 V_low
+ 3.267010000e-07 V_low
+ 3.268000000e-07 V_low
+ 3.268010000e-07 V_low
+ 3.269000000e-07 V_low
+ 3.269010000e-07 V_low
+ 3.270000000e-07 V_low
+ 3.270010000e-07 V_low
+ 3.271000000e-07 V_low
+ 3.271010000e-07 V_low
+ 3.272000000e-07 V_low
+ 3.272010000e-07 V_low
+ 3.273000000e-07 V_low
+ 3.273010000e-07 V_low
+ 3.274000000e-07 V_low
+ 3.274010000e-07 V_low
+ 3.275000000e-07 V_low
+ 3.275010000e-07 V_low
+ 3.276000000e-07 V_low
+ 3.276010000e-07 V_low
+ 3.277000000e-07 V_low
+ 3.277010000e-07 V_low
+ 3.278000000e-07 V_low
+ 3.278010000e-07 V_low
+ 3.279000000e-07 V_low
+ 3.279010000e-07 V_hig
+ 3.280000000e-07 V_hig
+ 3.280010000e-07 V_hig
+ 3.281000000e-07 V_hig
+ 3.281010000e-07 V_hig
+ 3.282000000e-07 V_hig
+ 3.282010000e-07 V_hig
+ 3.283000000e-07 V_hig
+ 3.283010000e-07 V_hig
+ 3.284000000e-07 V_hig
+ 3.284010000e-07 V_hig
+ 3.285000000e-07 V_hig
+ 3.285010000e-07 V_hig
+ 3.286000000e-07 V_hig
+ 3.286010000e-07 V_hig
+ 3.287000000e-07 V_hig
+ 3.287010000e-07 V_hig
+ 3.288000000e-07 V_hig
+ 3.288010000e-07 V_hig
+ 3.289000000e-07 V_hig
+ 3.289010000e-07 V_low
+ 3.290000000e-07 V_low
+ 3.290010000e-07 V_low
+ 3.291000000e-07 V_low
+ 3.291010000e-07 V_low
+ 3.292000000e-07 V_low
+ 3.292010000e-07 V_low
+ 3.293000000e-07 V_low
+ 3.293010000e-07 V_low
+ 3.294000000e-07 V_low
+ 3.294010000e-07 V_low
+ 3.295000000e-07 V_low
+ 3.295010000e-07 V_low
+ 3.296000000e-07 V_low
+ 3.296010000e-07 V_low
+ 3.297000000e-07 V_low
+ 3.297010000e-07 V_low
+ 3.298000000e-07 V_low
+ 3.298010000e-07 V_low
+ 3.299000000e-07 V_low
+ 3.299010000e-07 V_hig
+ 3.300000000e-07 V_hig
+ 3.300010000e-07 V_hig
+ 3.301000000e-07 V_hig
+ 3.301010000e-07 V_hig
+ 3.302000000e-07 V_hig
+ 3.302010000e-07 V_hig
+ 3.303000000e-07 V_hig
+ 3.303010000e-07 V_hig
+ 3.304000000e-07 V_hig
+ 3.304010000e-07 V_hig
+ 3.305000000e-07 V_hig
+ 3.305010000e-07 V_hig
+ 3.306000000e-07 V_hig
+ 3.306010000e-07 V_hig
+ 3.307000000e-07 V_hig
+ 3.307010000e-07 V_hig
+ 3.308000000e-07 V_hig
+ 3.308010000e-07 V_hig
+ 3.309000000e-07 V_hig
+ 3.309010000e-07 V_low
+ 3.310000000e-07 V_low
+ 3.310010000e-07 V_low
+ 3.311000000e-07 V_low
+ 3.311010000e-07 V_low
+ 3.312000000e-07 V_low
+ 3.312010000e-07 V_low
+ 3.313000000e-07 V_low
+ 3.313010000e-07 V_low
+ 3.314000000e-07 V_low
+ 3.314010000e-07 V_low
+ 3.315000000e-07 V_low
+ 3.315010000e-07 V_low
+ 3.316000000e-07 V_low
+ 3.316010000e-07 V_low
+ 3.317000000e-07 V_low
+ 3.317010000e-07 V_low
+ 3.318000000e-07 V_low
+ 3.318010000e-07 V_low
+ 3.319000000e-07 V_low
+ 3.319010000e-07 V_low
+ 3.320000000e-07 V_low
+ 3.320010000e-07 V_low
+ 3.321000000e-07 V_low
+ 3.321010000e-07 V_low
+ 3.322000000e-07 V_low
+ 3.322010000e-07 V_low
+ 3.323000000e-07 V_low
+ 3.323010000e-07 V_low
+ 3.324000000e-07 V_low
+ 3.324010000e-07 V_low
+ 3.325000000e-07 V_low
+ 3.325010000e-07 V_low
+ 3.326000000e-07 V_low
+ 3.326010000e-07 V_low
+ 3.327000000e-07 V_low
+ 3.327010000e-07 V_low
+ 3.328000000e-07 V_low
+ 3.328010000e-07 V_low
+ 3.329000000e-07 V_low
+ 3.329010000e-07 V_low
+ 3.330000000e-07 V_low
+ 3.330010000e-07 V_low
+ 3.331000000e-07 V_low
+ 3.331010000e-07 V_low
+ 3.332000000e-07 V_low
+ 3.332010000e-07 V_low
+ 3.333000000e-07 V_low
+ 3.333010000e-07 V_low
+ 3.334000000e-07 V_low
+ 3.334010000e-07 V_low
+ 3.335000000e-07 V_low
+ 3.335010000e-07 V_low
+ 3.336000000e-07 V_low
+ 3.336010000e-07 V_low
+ 3.337000000e-07 V_low
+ 3.337010000e-07 V_low
+ 3.338000000e-07 V_low
+ 3.338010000e-07 V_low
+ 3.339000000e-07 V_low
+ 3.339010000e-07 V_hig
+ 3.340000000e-07 V_hig
+ 3.340010000e-07 V_hig
+ 3.341000000e-07 V_hig
+ 3.341010000e-07 V_hig
+ 3.342000000e-07 V_hig
+ 3.342010000e-07 V_hig
+ 3.343000000e-07 V_hig
+ 3.343010000e-07 V_hig
+ 3.344000000e-07 V_hig
+ 3.344010000e-07 V_hig
+ 3.345000000e-07 V_hig
+ 3.345010000e-07 V_hig
+ 3.346000000e-07 V_hig
+ 3.346010000e-07 V_hig
+ 3.347000000e-07 V_hig
+ 3.347010000e-07 V_hig
+ 3.348000000e-07 V_hig
+ 3.348010000e-07 V_hig
+ 3.349000000e-07 V_hig
+ 3.349010000e-07 V_hig
+ 3.350000000e-07 V_hig
+ 3.350010000e-07 V_hig
+ 3.351000000e-07 V_hig
+ 3.351010000e-07 V_hig
+ 3.352000000e-07 V_hig
+ 3.352010000e-07 V_hig
+ 3.353000000e-07 V_hig
+ 3.353010000e-07 V_hig
+ 3.354000000e-07 V_hig
+ 3.354010000e-07 V_hig
+ 3.355000000e-07 V_hig
+ 3.355010000e-07 V_hig
+ 3.356000000e-07 V_hig
+ 3.356010000e-07 V_hig
+ 3.357000000e-07 V_hig
+ 3.357010000e-07 V_hig
+ 3.358000000e-07 V_hig
+ 3.358010000e-07 V_hig
+ 3.359000000e-07 V_hig
+ 3.359010000e-07 V_hig
+ 3.360000000e-07 V_hig
+ 3.360010000e-07 V_hig
+ 3.361000000e-07 V_hig
+ 3.361010000e-07 V_hig
+ 3.362000000e-07 V_hig
+ 3.362010000e-07 V_hig
+ 3.363000000e-07 V_hig
+ 3.363010000e-07 V_hig
+ 3.364000000e-07 V_hig
+ 3.364010000e-07 V_hig
+ 3.365000000e-07 V_hig
+ 3.365010000e-07 V_hig
+ 3.366000000e-07 V_hig
+ 3.366010000e-07 V_hig
+ 3.367000000e-07 V_hig
+ 3.367010000e-07 V_hig
+ 3.368000000e-07 V_hig
+ 3.368010000e-07 V_hig
+ 3.369000000e-07 V_hig
+ 3.369010000e-07 V_hig
+ 3.370000000e-07 V_hig
+ 3.370010000e-07 V_hig
+ 3.371000000e-07 V_hig
+ 3.371010000e-07 V_hig
+ 3.372000000e-07 V_hig
+ 3.372010000e-07 V_hig
+ 3.373000000e-07 V_hig
+ 3.373010000e-07 V_hig
+ 3.374000000e-07 V_hig
+ 3.374010000e-07 V_hig
+ 3.375000000e-07 V_hig
+ 3.375010000e-07 V_hig
+ 3.376000000e-07 V_hig
+ 3.376010000e-07 V_hig
+ 3.377000000e-07 V_hig
+ 3.377010000e-07 V_hig
+ 3.378000000e-07 V_hig
+ 3.378010000e-07 V_hig
+ 3.379000000e-07 V_hig
+ 3.379010000e-07 V_low
+ 3.380000000e-07 V_low
+ 3.380010000e-07 V_low
+ 3.381000000e-07 V_low
+ 3.381010000e-07 V_low
+ 3.382000000e-07 V_low
+ 3.382010000e-07 V_low
+ 3.383000000e-07 V_low
+ 3.383010000e-07 V_low
+ 3.384000000e-07 V_low
+ 3.384010000e-07 V_low
+ 3.385000000e-07 V_low
+ 3.385010000e-07 V_low
+ 3.386000000e-07 V_low
+ 3.386010000e-07 V_low
+ 3.387000000e-07 V_low
+ 3.387010000e-07 V_low
+ 3.388000000e-07 V_low
+ 3.388010000e-07 V_low
+ 3.389000000e-07 V_low
+ 3.389010000e-07 V_hig
+ 3.390000000e-07 V_hig
+ 3.390010000e-07 V_hig
+ 3.391000000e-07 V_hig
+ 3.391010000e-07 V_hig
+ 3.392000000e-07 V_hig
+ 3.392010000e-07 V_hig
+ 3.393000000e-07 V_hig
+ 3.393010000e-07 V_hig
+ 3.394000000e-07 V_hig
+ 3.394010000e-07 V_hig
+ 3.395000000e-07 V_hig
+ 3.395010000e-07 V_hig
+ 3.396000000e-07 V_hig
+ 3.396010000e-07 V_hig
+ 3.397000000e-07 V_hig
+ 3.397010000e-07 V_hig
+ 3.398000000e-07 V_hig
+ 3.398010000e-07 V_hig
+ 3.399000000e-07 V_hig
+ 3.399010000e-07 V_hig
+ 3.400000000e-07 V_hig
+ 3.400010000e-07 V_hig
+ 3.401000000e-07 V_hig
+ 3.401010000e-07 V_hig
+ 3.402000000e-07 V_hig
+ 3.402010000e-07 V_hig
+ 3.403000000e-07 V_hig
+ 3.403010000e-07 V_hig
+ 3.404000000e-07 V_hig
+ 3.404010000e-07 V_hig
+ 3.405000000e-07 V_hig
+ 3.405010000e-07 V_hig
+ 3.406000000e-07 V_hig
+ 3.406010000e-07 V_hig
+ 3.407000000e-07 V_hig
+ 3.407010000e-07 V_hig
+ 3.408000000e-07 V_hig
+ 3.408010000e-07 V_hig
+ 3.409000000e-07 V_hig
+ 3.409010000e-07 V_low
+ 3.410000000e-07 V_low
+ 3.410010000e-07 V_low
+ 3.411000000e-07 V_low
+ 3.411010000e-07 V_low
+ 3.412000000e-07 V_low
+ 3.412010000e-07 V_low
+ 3.413000000e-07 V_low
+ 3.413010000e-07 V_low
+ 3.414000000e-07 V_low
+ 3.414010000e-07 V_low
+ 3.415000000e-07 V_low
+ 3.415010000e-07 V_low
+ 3.416000000e-07 V_low
+ 3.416010000e-07 V_low
+ 3.417000000e-07 V_low
+ 3.417010000e-07 V_low
+ 3.418000000e-07 V_low
+ 3.418010000e-07 V_low
+ 3.419000000e-07 V_low
+ 3.419010000e-07 V_hig
+ 3.420000000e-07 V_hig
+ 3.420010000e-07 V_hig
+ 3.421000000e-07 V_hig
+ 3.421010000e-07 V_hig
+ 3.422000000e-07 V_hig
+ 3.422010000e-07 V_hig
+ 3.423000000e-07 V_hig
+ 3.423010000e-07 V_hig
+ 3.424000000e-07 V_hig
+ 3.424010000e-07 V_hig
+ 3.425000000e-07 V_hig
+ 3.425010000e-07 V_hig
+ 3.426000000e-07 V_hig
+ 3.426010000e-07 V_hig
+ 3.427000000e-07 V_hig
+ 3.427010000e-07 V_hig
+ 3.428000000e-07 V_hig
+ 3.428010000e-07 V_hig
+ 3.429000000e-07 V_hig
+ 3.429010000e-07 V_hig
+ 3.430000000e-07 V_hig
+ 3.430010000e-07 V_hig
+ 3.431000000e-07 V_hig
+ 3.431010000e-07 V_hig
+ 3.432000000e-07 V_hig
+ 3.432010000e-07 V_hig
+ 3.433000000e-07 V_hig
+ 3.433010000e-07 V_hig
+ 3.434000000e-07 V_hig
+ 3.434010000e-07 V_hig
+ 3.435000000e-07 V_hig
+ 3.435010000e-07 V_hig
+ 3.436000000e-07 V_hig
+ 3.436010000e-07 V_hig
+ 3.437000000e-07 V_hig
+ 3.437010000e-07 V_hig
+ 3.438000000e-07 V_hig
+ 3.438010000e-07 V_hig
+ 3.439000000e-07 V_hig
+ 3.439010000e-07 V_hig
+ 3.440000000e-07 V_hig
+ 3.440010000e-07 V_hig
+ 3.441000000e-07 V_hig
+ 3.441010000e-07 V_hig
+ 3.442000000e-07 V_hig
+ 3.442010000e-07 V_hig
+ 3.443000000e-07 V_hig
+ 3.443010000e-07 V_hig
+ 3.444000000e-07 V_hig
+ 3.444010000e-07 V_hig
+ 3.445000000e-07 V_hig
+ 3.445010000e-07 V_hig
+ 3.446000000e-07 V_hig
+ 3.446010000e-07 V_hig
+ 3.447000000e-07 V_hig
+ 3.447010000e-07 V_hig
+ 3.448000000e-07 V_hig
+ 3.448010000e-07 V_hig
+ 3.449000000e-07 V_hig
+ 3.449010000e-07 V_hig
+ 3.450000000e-07 V_hig
+ 3.450010000e-07 V_hig
+ 3.451000000e-07 V_hig
+ 3.451010000e-07 V_hig
+ 3.452000000e-07 V_hig
+ 3.452010000e-07 V_hig
+ 3.453000000e-07 V_hig
+ 3.453010000e-07 V_hig
+ 3.454000000e-07 V_hig
+ 3.454010000e-07 V_hig
+ 3.455000000e-07 V_hig
+ 3.455010000e-07 V_hig
+ 3.456000000e-07 V_hig
+ 3.456010000e-07 V_hig
+ 3.457000000e-07 V_hig
+ 3.457010000e-07 V_hig
+ 3.458000000e-07 V_hig
+ 3.458010000e-07 V_hig
+ 3.459000000e-07 V_hig
+ 3.459010000e-07 V_low
+ 3.460000000e-07 V_low
+ 3.460010000e-07 V_low
+ 3.461000000e-07 V_low
+ 3.461010000e-07 V_low
+ 3.462000000e-07 V_low
+ 3.462010000e-07 V_low
+ 3.463000000e-07 V_low
+ 3.463010000e-07 V_low
+ 3.464000000e-07 V_low
+ 3.464010000e-07 V_low
+ 3.465000000e-07 V_low
+ 3.465010000e-07 V_low
+ 3.466000000e-07 V_low
+ 3.466010000e-07 V_low
+ 3.467000000e-07 V_low
+ 3.467010000e-07 V_low
+ 3.468000000e-07 V_low
+ 3.468010000e-07 V_low
+ 3.469000000e-07 V_low
+ 3.469010000e-07 V_low
+ 3.470000000e-07 V_low
+ 3.470010000e-07 V_low
+ 3.471000000e-07 V_low
+ 3.471010000e-07 V_low
+ 3.472000000e-07 V_low
+ 3.472010000e-07 V_low
+ 3.473000000e-07 V_low
+ 3.473010000e-07 V_low
+ 3.474000000e-07 V_low
+ 3.474010000e-07 V_low
+ 3.475000000e-07 V_low
+ 3.475010000e-07 V_low
+ 3.476000000e-07 V_low
+ 3.476010000e-07 V_low
+ 3.477000000e-07 V_low
+ 3.477010000e-07 V_low
+ 3.478000000e-07 V_low
+ 3.478010000e-07 V_low
+ 3.479000000e-07 V_low
+ 3.479010000e-07 V_low
+ 3.480000000e-07 V_low
+ 3.480010000e-07 V_low
+ 3.481000000e-07 V_low
+ 3.481010000e-07 V_low
+ 3.482000000e-07 V_low
+ 3.482010000e-07 V_low
+ 3.483000000e-07 V_low
+ 3.483010000e-07 V_low
+ 3.484000000e-07 V_low
+ 3.484010000e-07 V_low
+ 3.485000000e-07 V_low
+ 3.485010000e-07 V_low
+ 3.486000000e-07 V_low
+ 3.486010000e-07 V_low
+ 3.487000000e-07 V_low
+ 3.487010000e-07 V_low
+ 3.488000000e-07 V_low
+ 3.488010000e-07 V_low
+ 3.489000000e-07 V_low
+ 3.489010000e-07 V_low
+ 3.490000000e-07 V_low
+ 3.490010000e-07 V_low
+ 3.491000000e-07 V_low
+ 3.491010000e-07 V_low
+ 3.492000000e-07 V_low
+ 3.492010000e-07 V_low
+ 3.493000000e-07 V_low
+ 3.493010000e-07 V_low
+ 3.494000000e-07 V_low
+ 3.494010000e-07 V_low
+ 3.495000000e-07 V_low
+ 3.495010000e-07 V_low
+ 3.496000000e-07 V_low
+ 3.496010000e-07 V_low
+ 3.497000000e-07 V_low
+ 3.497010000e-07 V_low
+ 3.498000000e-07 V_low
+ 3.498010000e-07 V_low
+ 3.499000000e-07 V_low
+ 3.499010000e-07 V_low
+ 3.500000000e-07 V_low
+ 3.500010000e-07 V_low
+ 3.501000000e-07 V_low
+ 3.501010000e-07 V_low
+ 3.502000000e-07 V_low
+ 3.502010000e-07 V_low
+ 3.503000000e-07 V_low
+ 3.503010000e-07 V_low
+ 3.504000000e-07 V_low
+ 3.504010000e-07 V_low
+ 3.505000000e-07 V_low
+ 3.505010000e-07 V_low
+ 3.506000000e-07 V_low
+ 3.506010000e-07 V_low
+ 3.507000000e-07 V_low
+ 3.507010000e-07 V_low
+ 3.508000000e-07 V_low
+ 3.508010000e-07 V_low
+ 3.509000000e-07 V_low
+ 3.509010000e-07 V_hig
+ 3.510000000e-07 V_hig
+ 3.510010000e-07 V_hig
+ 3.511000000e-07 V_hig
+ 3.511010000e-07 V_hig
+ 3.512000000e-07 V_hig
+ 3.512010000e-07 V_hig
+ 3.513000000e-07 V_hig
+ 3.513010000e-07 V_hig
+ 3.514000000e-07 V_hig
+ 3.514010000e-07 V_hig
+ 3.515000000e-07 V_hig
+ 3.515010000e-07 V_hig
+ 3.516000000e-07 V_hig
+ 3.516010000e-07 V_hig
+ 3.517000000e-07 V_hig
+ 3.517010000e-07 V_hig
+ 3.518000000e-07 V_hig
+ 3.518010000e-07 V_hig
+ 3.519000000e-07 V_hig
+ 3.519010000e-07 V_hig
+ 3.520000000e-07 V_hig
+ 3.520010000e-07 V_hig
+ 3.521000000e-07 V_hig
+ 3.521010000e-07 V_hig
+ 3.522000000e-07 V_hig
+ 3.522010000e-07 V_hig
+ 3.523000000e-07 V_hig
+ 3.523010000e-07 V_hig
+ 3.524000000e-07 V_hig
+ 3.524010000e-07 V_hig
+ 3.525000000e-07 V_hig
+ 3.525010000e-07 V_hig
+ 3.526000000e-07 V_hig
+ 3.526010000e-07 V_hig
+ 3.527000000e-07 V_hig
+ 3.527010000e-07 V_hig
+ 3.528000000e-07 V_hig
+ 3.528010000e-07 V_hig
+ 3.529000000e-07 V_hig
+ 3.529010000e-07 V_low
+ 3.530000000e-07 V_low
+ 3.530010000e-07 V_low
+ 3.531000000e-07 V_low
+ 3.531010000e-07 V_low
+ 3.532000000e-07 V_low
+ 3.532010000e-07 V_low
+ 3.533000000e-07 V_low
+ 3.533010000e-07 V_low
+ 3.534000000e-07 V_low
+ 3.534010000e-07 V_low
+ 3.535000000e-07 V_low
+ 3.535010000e-07 V_low
+ 3.536000000e-07 V_low
+ 3.536010000e-07 V_low
+ 3.537000000e-07 V_low
+ 3.537010000e-07 V_low
+ 3.538000000e-07 V_low
+ 3.538010000e-07 V_low
+ 3.539000000e-07 V_low
+ 3.539010000e-07 V_hig
+ 3.540000000e-07 V_hig
+ 3.540010000e-07 V_hig
+ 3.541000000e-07 V_hig
+ 3.541010000e-07 V_hig
+ 3.542000000e-07 V_hig
+ 3.542010000e-07 V_hig
+ 3.543000000e-07 V_hig
+ 3.543010000e-07 V_hig
+ 3.544000000e-07 V_hig
+ 3.544010000e-07 V_hig
+ 3.545000000e-07 V_hig
+ 3.545010000e-07 V_hig
+ 3.546000000e-07 V_hig
+ 3.546010000e-07 V_hig
+ 3.547000000e-07 V_hig
+ 3.547010000e-07 V_hig
+ 3.548000000e-07 V_hig
+ 3.548010000e-07 V_hig
+ 3.549000000e-07 V_hig
+ 3.549010000e-07 V_hig
+ 3.550000000e-07 V_hig
+ 3.550010000e-07 V_hig
+ 3.551000000e-07 V_hig
+ 3.551010000e-07 V_hig
+ 3.552000000e-07 V_hig
+ 3.552010000e-07 V_hig
+ 3.553000000e-07 V_hig
+ 3.553010000e-07 V_hig
+ 3.554000000e-07 V_hig
+ 3.554010000e-07 V_hig
+ 3.555000000e-07 V_hig
+ 3.555010000e-07 V_hig
+ 3.556000000e-07 V_hig
+ 3.556010000e-07 V_hig
+ 3.557000000e-07 V_hig
+ 3.557010000e-07 V_hig
+ 3.558000000e-07 V_hig
+ 3.558010000e-07 V_hig
+ 3.559000000e-07 V_hig
+ 3.559010000e-07 V_low
+ 3.560000000e-07 V_low
+ 3.560010000e-07 V_low
+ 3.561000000e-07 V_low
+ 3.561010000e-07 V_low
+ 3.562000000e-07 V_low
+ 3.562010000e-07 V_low
+ 3.563000000e-07 V_low
+ 3.563010000e-07 V_low
+ 3.564000000e-07 V_low
+ 3.564010000e-07 V_low
+ 3.565000000e-07 V_low
+ 3.565010000e-07 V_low
+ 3.566000000e-07 V_low
+ 3.566010000e-07 V_low
+ 3.567000000e-07 V_low
+ 3.567010000e-07 V_low
+ 3.568000000e-07 V_low
+ 3.568010000e-07 V_low
+ 3.569000000e-07 V_low
+ 3.569010000e-07 V_low
+ 3.570000000e-07 V_low
+ 3.570010000e-07 V_low
+ 3.571000000e-07 V_low
+ 3.571010000e-07 V_low
+ 3.572000000e-07 V_low
+ 3.572010000e-07 V_low
+ 3.573000000e-07 V_low
+ 3.573010000e-07 V_low
+ 3.574000000e-07 V_low
+ 3.574010000e-07 V_low
+ 3.575000000e-07 V_low
+ 3.575010000e-07 V_low
+ 3.576000000e-07 V_low
+ 3.576010000e-07 V_low
+ 3.577000000e-07 V_low
+ 3.577010000e-07 V_low
+ 3.578000000e-07 V_low
+ 3.578010000e-07 V_low
+ 3.579000000e-07 V_low
+ 3.579010000e-07 V_low
+ 3.580000000e-07 V_low
+ 3.580010000e-07 V_low
+ 3.581000000e-07 V_low
+ 3.581010000e-07 V_low
+ 3.582000000e-07 V_low
+ 3.582010000e-07 V_low
+ 3.583000000e-07 V_low
+ 3.583010000e-07 V_low
+ 3.584000000e-07 V_low
+ 3.584010000e-07 V_low
+ 3.585000000e-07 V_low
+ 3.585010000e-07 V_low
+ 3.586000000e-07 V_low
+ 3.586010000e-07 V_low
+ 3.587000000e-07 V_low
+ 3.587010000e-07 V_low
+ 3.588000000e-07 V_low
+ 3.588010000e-07 V_low
+ 3.589000000e-07 V_low
+ 3.589010000e-07 V_low
+ 3.590000000e-07 V_low
+ 3.590010000e-07 V_low
+ 3.591000000e-07 V_low
+ 3.591010000e-07 V_low
+ 3.592000000e-07 V_low
+ 3.592010000e-07 V_low
+ 3.593000000e-07 V_low
+ 3.593010000e-07 V_low
+ 3.594000000e-07 V_low
+ 3.594010000e-07 V_low
+ 3.595000000e-07 V_low
+ 3.595010000e-07 V_low
+ 3.596000000e-07 V_low
+ 3.596010000e-07 V_low
+ 3.597000000e-07 V_low
+ 3.597010000e-07 V_low
+ 3.598000000e-07 V_low
+ 3.598010000e-07 V_low
+ 3.599000000e-07 V_low
+ 3.599010000e-07 V_hig
+ 3.600000000e-07 V_hig
+ 3.600010000e-07 V_hig
+ 3.601000000e-07 V_hig
+ 3.601010000e-07 V_hig
+ 3.602000000e-07 V_hig
+ 3.602010000e-07 V_hig
+ 3.603000000e-07 V_hig
+ 3.603010000e-07 V_hig
+ 3.604000000e-07 V_hig
+ 3.604010000e-07 V_hig
+ 3.605000000e-07 V_hig
+ 3.605010000e-07 V_hig
+ 3.606000000e-07 V_hig
+ 3.606010000e-07 V_hig
+ 3.607000000e-07 V_hig
+ 3.607010000e-07 V_hig
+ 3.608000000e-07 V_hig
+ 3.608010000e-07 V_hig
+ 3.609000000e-07 V_hig
+ 3.609010000e-07 V_low
+ 3.610000000e-07 V_low
+ 3.610010000e-07 V_low
+ 3.611000000e-07 V_low
+ 3.611010000e-07 V_low
+ 3.612000000e-07 V_low
+ 3.612010000e-07 V_low
+ 3.613000000e-07 V_low
+ 3.613010000e-07 V_low
+ 3.614000000e-07 V_low
+ 3.614010000e-07 V_low
+ 3.615000000e-07 V_low
+ 3.615010000e-07 V_low
+ 3.616000000e-07 V_low
+ 3.616010000e-07 V_low
+ 3.617000000e-07 V_low
+ 3.617010000e-07 V_low
+ 3.618000000e-07 V_low
+ 3.618010000e-07 V_low
+ 3.619000000e-07 V_low
+ 3.619010000e-07 V_hig
+ 3.620000000e-07 V_hig
+ 3.620010000e-07 V_hig
+ 3.621000000e-07 V_hig
+ 3.621010000e-07 V_hig
+ 3.622000000e-07 V_hig
+ 3.622010000e-07 V_hig
+ 3.623000000e-07 V_hig
+ 3.623010000e-07 V_hig
+ 3.624000000e-07 V_hig
+ 3.624010000e-07 V_hig
+ 3.625000000e-07 V_hig
+ 3.625010000e-07 V_hig
+ 3.626000000e-07 V_hig
+ 3.626010000e-07 V_hig
+ 3.627000000e-07 V_hig
+ 3.627010000e-07 V_hig
+ 3.628000000e-07 V_hig
+ 3.628010000e-07 V_hig
+ 3.629000000e-07 V_hig
+ 3.629010000e-07 V_hig
+ 3.630000000e-07 V_hig
+ 3.630010000e-07 V_hig
+ 3.631000000e-07 V_hig
+ 3.631010000e-07 V_hig
+ 3.632000000e-07 V_hig
+ 3.632010000e-07 V_hig
+ 3.633000000e-07 V_hig
+ 3.633010000e-07 V_hig
+ 3.634000000e-07 V_hig
+ 3.634010000e-07 V_hig
+ 3.635000000e-07 V_hig
+ 3.635010000e-07 V_hig
+ 3.636000000e-07 V_hig
+ 3.636010000e-07 V_hig
+ 3.637000000e-07 V_hig
+ 3.637010000e-07 V_hig
+ 3.638000000e-07 V_hig
+ 3.638010000e-07 V_hig
+ 3.639000000e-07 V_hig
+ 3.639010000e-07 V_low
+ 3.640000000e-07 V_low
+ 3.640010000e-07 V_low
+ 3.641000000e-07 V_low
+ 3.641010000e-07 V_low
+ 3.642000000e-07 V_low
+ 3.642010000e-07 V_low
+ 3.643000000e-07 V_low
+ 3.643010000e-07 V_low
+ 3.644000000e-07 V_low
+ 3.644010000e-07 V_low
+ 3.645000000e-07 V_low
+ 3.645010000e-07 V_low
+ 3.646000000e-07 V_low
+ 3.646010000e-07 V_low
+ 3.647000000e-07 V_low
+ 3.647010000e-07 V_low
+ 3.648000000e-07 V_low
+ 3.648010000e-07 V_low
+ 3.649000000e-07 V_low
+ 3.649010000e-07 V_hig
+ 3.650000000e-07 V_hig
+ 3.650010000e-07 V_hig
+ 3.651000000e-07 V_hig
+ 3.651010000e-07 V_hig
+ 3.652000000e-07 V_hig
+ 3.652010000e-07 V_hig
+ 3.653000000e-07 V_hig
+ 3.653010000e-07 V_hig
+ 3.654000000e-07 V_hig
+ 3.654010000e-07 V_hig
+ 3.655000000e-07 V_hig
+ 3.655010000e-07 V_hig
+ 3.656000000e-07 V_hig
+ 3.656010000e-07 V_hig
+ 3.657000000e-07 V_hig
+ 3.657010000e-07 V_hig
+ 3.658000000e-07 V_hig
+ 3.658010000e-07 V_hig
+ 3.659000000e-07 V_hig
+ 3.659010000e-07 V_low
+ 3.660000000e-07 V_low
+ 3.660010000e-07 V_low
+ 3.661000000e-07 V_low
+ 3.661010000e-07 V_low
+ 3.662000000e-07 V_low
+ 3.662010000e-07 V_low
+ 3.663000000e-07 V_low
+ 3.663010000e-07 V_low
+ 3.664000000e-07 V_low
+ 3.664010000e-07 V_low
+ 3.665000000e-07 V_low
+ 3.665010000e-07 V_low
+ 3.666000000e-07 V_low
+ 3.666010000e-07 V_low
+ 3.667000000e-07 V_low
+ 3.667010000e-07 V_low
+ 3.668000000e-07 V_low
+ 3.668010000e-07 V_low
+ 3.669000000e-07 V_low
+ 3.669010000e-07 V_low
+ 3.670000000e-07 V_low
+ 3.670010000e-07 V_low
+ 3.671000000e-07 V_low
+ 3.671010000e-07 V_low
+ 3.672000000e-07 V_low
+ 3.672010000e-07 V_low
+ 3.673000000e-07 V_low
+ 3.673010000e-07 V_low
+ 3.674000000e-07 V_low
+ 3.674010000e-07 V_low
+ 3.675000000e-07 V_low
+ 3.675010000e-07 V_low
+ 3.676000000e-07 V_low
+ 3.676010000e-07 V_low
+ 3.677000000e-07 V_low
+ 3.677010000e-07 V_low
+ 3.678000000e-07 V_low
+ 3.678010000e-07 V_low
+ 3.679000000e-07 V_low
+ 3.679010000e-07 V_low
+ 3.680000000e-07 V_low
+ 3.680010000e-07 V_low
+ 3.681000000e-07 V_low
+ 3.681010000e-07 V_low
+ 3.682000000e-07 V_low
+ 3.682010000e-07 V_low
+ 3.683000000e-07 V_low
+ 3.683010000e-07 V_low
+ 3.684000000e-07 V_low
+ 3.684010000e-07 V_low
+ 3.685000000e-07 V_low
+ 3.685010000e-07 V_low
+ 3.686000000e-07 V_low
+ 3.686010000e-07 V_low
+ 3.687000000e-07 V_low
+ 3.687010000e-07 V_low
+ 3.688000000e-07 V_low
+ 3.688010000e-07 V_low
+ 3.689000000e-07 V_low
+ 3.689010000e-07 V_hig
+ 3.690000000e-07 V_hig
+ 3.690010000e-07 V_hig
+ 3.691000000e-07 V_hig
+ 3.691010000e-07 V_hig
+ 3.692000000e-07 V_hig
+ 3.692010000e-07 V_hig
+ 3.693000000e-07 V_hig
+ 3.693010000e-07 V_hig
+ 3.694000000e-07 V_hig
+ 3.694010000e-07 V_hig
+ 3.695000000e-07 V_hig
+ 3.695010000e-07 V_hig
+ 3.696000000e-07 V_hig
+ 3.696010000e-07 V_hig
+ 3.697000000e-07 V_hig
+ 3.697010000e-07 V_hig
+ 3.698000000e-07 V_hig
+ 3.698010000e-07 V_hig
+ 3.699000000e-07 V_hig
+ 3.699010000e-07 V_hig
+ 3.700000000e-07 V_hig
+ 3.700010000e-07 V_hig
+ 3.701000000e-07 V_hig
+ 3.701010000e-07 V_hig
+ 3.702000000e-07 V_hig
+ 3.702010000e-07 V_hig
+ 3.703000000e-07 V_hig
+ 3.703010000e-07 V_hig
+ 3.704000000e-07 V_hig
+ 3.704010000e-07 V_hig
+ 3.705000000e-07 V_hig
+ 3.705010000e-07 V_hig
+ 3.706000000e-07 V_hig
+ 3.706010000e-07 V_hig
+ 3.707000000e-07 V_hig
+ 3.707010000e-07 V_hig
+ 3.708000000e-07 V_hig
+ 3.708010000e-07 V_hig
+ 3.709000000e-07 V_hig
+ 3.709010000e-07 V_low
+ 3.710000000e-07 V_low
+ 3.710010000e-07 V_low
+ 3.711000000e-07 V_low
+ 3.711010000e-07 V_low
+ 3.712000000e-07 V_low
+ 3.712010000e-07 V_low
+ 3.713000000e-07 V_low
+ 3.713010000e-07 V_low
+ 3.714000000e-07 V_low
+ 3.714010000e-07 V_low
+ 3.715000000e-07 V_low
+ 3.715010000e-07 V_low
+ 3.716000000e-07 V_low
+ 3.716010000e-07 V_low
+ 3.717000000e-07 V_low
+ 3.717010000e-07 V_low
+ 3.718000000e-07 V_low
+ 3.718010000e-07 V_low
+ 3.719000000e-07 V_low
+ 3.719010000e-07 V_low
+ 3.720000000e-07 V_low
+ 3.720010000e-07 V_low
+ 3.721000000e-07 V_low
+ 3.721010000e-07 V_low
+ 3.722000000e-07 V_low
+ 3.722010000e-07 V_low
+ 3.723000000e-07 V_low
+ 3.723010000e-07 V_low
+ 3.724000000e-07 V_low
+ 3.724010000e-07 V_low
+ 3.725000000e-07 V_low
+ 3.725010000e-07 V_low
+ 3.726000000e-07 V_low
+ 3.726010000e-07 V_low
+ 3.727000000e-07 V_low
+ 3.727010000e-07 V_low
+ 3.728000000e-07 V_low
+ 3.728010000e-07 V_low
+ 3.729000000e-07 V_low
+ 3.729010000e-07 V_hig
+ 3.730000000e-07 V_hig
+ 3.730010000e-07 V_hig
+ 3.731000000e-07 V_hig
+ 3.731010000e-07 V_hig
+ 3.732000000e-07 V_hig
+ 3.732010000e-07 V_hig
+ 3.733000000e-07 V_hig
+ 3.733010000e-07 V_hig
+ 3.734000000e-07 V_hig
+ 3.734010000e-07 V_hig
+ 3.735000000e-07 V_hig
+ 3.735010000e-07 V_hig
+ 3.736000000e-07 V_hig
+ 3.736010000e-07 V_hig
+ 3.737000000e-07 V_hig
+ 3.737010000e-07 V_hig
+ 3.738000000e-07 V_hig
+ 3.738010000e-07 V_hig
+ 3.739000000e-07 V_hig
+ 3.739010000e-07 V_low
+ 3.740000000e-07 V_low
+ 3.740010000e-07 V_low
+ 3.741000000e-07 V_low
+ 3.741010000e-07 V_low
+ 3.742000000e-07 V_low
+ 3.742010000e-07 V_low
+ 3.743000000e-07 V_low
+ 3.743010000e-07 V_low
+ 3.744000000e-07 V_low
+ 3.744010000e-07 V_low
+ 3.745000000e-07 V_low
+ 3.745010000e-07 V_low
+ 3.746000000e-07 V_low
+ 3.746010000e-07 V_low
+ 3.747000000e-07 V_low
+ 3.747010000e-07 V_low
+ 3.748000000e-07 V_low
+ 3.748010000e-07 V_low
+ 3.749000000e-07 V_low
+ 3.749010000e-07 V_low
+ 3.750000000e-07 V_low
+ 3.750010000e-07 V_low
+ 3.751000000e-07 V_low
+ 3.751010000e-07 V_low
+ 3.752000000e-07 V_low
+ 3.752010000e-07 V_low
+ 3.753000000e-07 V_low
+ 3.753010000e-07 V_low
+ 3.754000000e-07 V_low
+ 3.754010000e-07 V_low
+ 3.755000000e-07 V_low
+ 3.755010000e-07 V_low
+ 3.756000000e-07 V_low
+ 3.756010000e-07 V_low
+ 3.757000000e-07 V_low
+ 3.757010000e-07 V_low
+ 3.758000000e-07 V_low
+ 3.758010000e-07 V_low
+ 3.759000000e-07 V_low
+ 3.759010000e-07 V_hig
+ 3.760000000e-07 V_hig
+ 3.760010000e-07 V_hig
+ 3.761000000e-07 V_hig
+ 3.761010000e-07 V_hig
+ 3.762000000e-07 V_hig
+ 3.762010000e-07 V_hig
+ 3.763000000e-07 V_hig
+ 3.763010000e-07 V_hig
+ 3.764000000e-07 V_hig
+ 3.764010000e-07 V_hig
+ 3.765000000e-07 V_hig
+ 3.765010000e-07 V_hig
+ 3.766000000e-07 V_hig
+ 3.766010000e-07 V_hig
+ 3.767000000e-07 V_hig
+ 3.767010000e-07 V_hig
+ 3.768000000e-07 V_hig
+ 3.768010000e-07 V_hig
+ 3.769000000e-07 V_hig
+ 3.769010000e-07 V_hig
+ 3.770000000e-07 V_hig
+ 3.770010000e-07 V_hig
+ 3.771000000e-07 V_hig
+ 3.771010000e-07 V_hig
+ 3.772000000e-07 V_hig
+ 3.772010000e-07 V_hig
+ 3.773000000e-07 V_hig
+ 3.773010000e-07 V_hig
+ 3.774000000e-07 V_hig
+ 3.774010000e-07 V_hig
+ 3.775000000e-07 V_hig
+ 3.775010000e-07 V_hig
+ 3.776000000e-07 V_hig
+ 3.776010000e-07 V_hig
+ 3.777000000e-07 V_hig
+ 3.777010000e-07 V_hig
+ 3.778000000e-07 V_hig
+ 3.778010000e-07 V_hig
+ 3.779000000e-07 V_hig
+ 3.779010000e-07 V_low
+ 3.780000000e-07 V_low
+ 3.780010000e-07 V_low
+ 3.781000000e-07 V_low
+ 3.781010000e-07 V_low
+ 3.782000000e-07 V_low
+ 3.782010000e-07 V_low
+ 3.783000000e-07 V_low
+ 3.783010000e-07 V_low
+ 3.784000000e-07 V_low
+ 3.784010000e-07 V_low
+ 3.785000000e-07 V_low
+ 3.785010000e-07 V_low
+ 3.786000000e-07 V_low
+ 3.786010000e-07 V_low
+ 3.787000000e-07 V_low
+ 3.787010000e-07 V_low
+ 3.788000000e-07 V_low
+ 3.788010000e-07 V_low
+ 3.789000000e-07 V_low
+ 3.789010000e-07 V_hig
+ 3.790000000e-07 V_hig
+ 3.790010000e-07 V_hig
+ 3.791000000e-07 V_hig
+ 3.791010000e-07 V_hig
+ 3.792000000e-07 V_hig
+ 3.792010000e-07 V_hig
+ 3.793000000e-07 V_hig
+ 3.793010000e-07 V_hig
+ 3.794000000e-07 V_hig
+ 3.794010000e-07 V_hig
+ 3.795000000e-07 V_hig
+ 3.795010000e-07 V_hig
+ 3.796000000e-07 V_hig
+ 3.796010000e-07 V_hig
+ 3.797000000e-07 V_hig
+ 3.797010000e-07 V_hig
+ 3.798000000e-07 V_hig
+ 3.798010000e-07 V_hig
+ 3.799000000e-07 V_hig
+ 3.799010000e-07 V_low
+ 3.800000000e-07 V_low
+ 3.800010000e-07 V_low
+ 3.801000000e-07 V_low
+ 3.801010000e-07 V_low
+ 3.802000000e-07 V_low
+ 3.802010000e-07 V_low
+ 3.803000000e-07 V_low
+ 3.803010000e-07 V_low
+ 3.804000000e-07 V_low
+ 3.804010000e-07 V_low
+ 3.805000000e-07 V_low
+ 3.805010000e-07 V_low
+ 3.806000000e-07 V_low
+ 3.806010000e-07 V_low
+ 3.807000000e-07 V_low
+ 3.807010000e-07 V_low
+ 3.808000000e-07 V_low
+ 3.808010000e-07 V_low
+ 3.809000000e-07 V_low
+ 3.809010000e-07 V_low
+ 3.810000000e-07 V_low
+ 3.810010000e-07 V_low
+ 3.811000000e-07 V_low
+ 3.811010000e-07 V_low
+ 3.812000000e-07 V_low
+ 3.812010000e-07 V_low
+ 3.813000000e-07 V_low
+ 3.813010000e-07 V_low
+ 3.814000000e-07 V_low
+ 3.814010000e-07 V_low
+ 3.815000000e-07 V_low
+ 3.815010000e-07 V_low
+ 3.816000000e-07 V_low
+ 3.816010000e-07 V_low
+ 3.817000000e-07 V_low
+ 3.817010000e-07 V_low
+ 3.818000000e-07 V_low
+ 3.818010000e-07 V_low
+ 3.819000000e-07 V_low
+ 3.819010000e-07 V_hig
+ 3.820000000e-07 V_hig
+ 3.820010000e-07 V_hig
+ 3.821000000e-07 V_hig
+ 3.821010000e-07 V_hig
+ 3.822000000e-07 V_hig
+ 3.822010000e-07 V_hig
+ 3.823000000e-07 V_hig
+ 3.823010000e-07 V_hig
+ 3.824000000e-07 V_hig
+ 3.824010000e-07 V_hig
+ 3.825000000e-07 V_hig
+ 3.825010000e-07 V_hig
+ 3.826000000e-07 V_hig
+ 3.826010000e-07 V_hig
+ 3.827000000e-07 V_hig
+ 3.827010000e-07 V_hig
+ 3.828000000e-07 V_hig
+ 3.828010000e-07 V_hig
+ 3.829000000e-07 V_hig
+ 3.829010000e-07 V_low
+ 3.830000000e-07 V_low
+ 3.830010000e-07 V_low
+ 3.831000000e-07 V_low
+ 3.831010000e-07 V_low
+ 3.832000000e-07 V_low
+ 3.832010000e-07 V_low
+ 3.833000000e-07 V_low
+ 3.833010000e-07 V_low
+ 3.834000000e-07 V_low
+ 3.834010000e-07 V_low
+ 3.835000000e-07 V_low
+ 3.835010000e-07 V_low
+ 3.836000000e-07 V_low
+ 3.836010000e-07 V_low
+ 3.837000000e-07 V_low
+ 3.837010000e-07 V_low
+ 3.838000000e-07 V_low
+ 3.838010000e-07 V_low
+ 3.839000000e-07 V_low
+ 3.839010000e-07 V_hig
+ 3.840000000e-07 V_hig
+ 3.840010000e-07 V_hig
+ 3.841000000e-07 V_hig
+ 3.841010000e-07 V_hig
+ 3.842000000e-07 V_hig
+ 3.842010000e-07 V_hig
+ 3.843000000e-07 V_hig
+ 3.843010000e-07 V_hig
+ 3.844000000e-07 V_hig
+ 3.844010000e-07 V_hig
+ 3.845000000e-07 V_hig
+ 3.845010000e-07 V_hig
+ 3.846000000e-07 V_hig
+ 3.846010000e-07 V_hig
+ 3.847000000e-07 V_hig
+ 3.847010000e-07 V_hig
+ 3.848000000e-07 V_hig
+ 3.848010000e-07 V_hig
+ 3.849000000e-07 V_hig
+ 3.849010000e-07 V_hig
+ 3.850000000e-07 V_hig
+ 3.850010000e-07 V_hig
+ 3.851000000e-07 V_hig
+ 3.851010000e-07 V_hig
+ 3.852000000e-07 V_hig
+ 3.852010000e-07 V_hig
+ 3.853000000e-07 V_hig
+ 3.853010000e-07 V_hig
+ 3.854000000e-07 V_hig
+ 3.854010000e-07 V_hig
+ 3.855000000e-07 V_hig
+ 3.855010000e-07 V_hig
+ 3.856000000e-07 V_hig
+ 3.856010000e-07 V_hig
+ 3.857000000e-07 V_hig
+ 3.857010000e-07 V_hig
+ 3.858000000e-07 V_hig
+ 3.858010000e-07 V_hig
+ 3.859000000e-07 V_hig
+ 3.859010000e-07 V_hig
+ 3.860000000e-07 V_hig
+ 3.860010000e-07 V_hig
+ 3.861000000e-07 V_hig
+ 3.861010000e-07 V_hig
+ 3.862000000e-07 V_hig
+ 3.862010000e-07 V_hig
+ 3.863000000e-07 V_hig
+ 3.863010000e-07 V_hig
+ 3.864000000e-07 V_hig
+ 3.864010000e-07 V_hig
+ 3.865000000e-07 V_hig
+ 3.865010000e-07 V_hig
+ 3.866000000e-07 V_hig
+ 3.866010000e-07 V_hig
+ 3.867000000e-07 V_hig
+ 3.867010000e-07 V_hig
+ 3.868000000e-07 V_hig
+ 3.868010000e-07 V_hig
+ 3.869000000e-07 V_hig
+ 3.869010000e-07 V_hig
+ 3.870000000e-07 V_hig
+ 3.870010000e-07 V_hig
+ 3.871000000e-07 V_hig
+ 3.871010000e-07 V_hig
+ 3.872000000e-07 V_hig
+ 3.872010000e-07 V_hig
+ 3.873000000e-07 V_hig
+ 3.873010000e-07 V_hig
+ 3.874000000e-07 V_hig
+ 3.874010000e-07 V_hig
+ 3.875000000e-07 V_hig
+ 3.875010000e-07 V_hig
+ 3.876000000e-07 V_hig
+ 3.876010000e-07 V_hig
+ 3.877000000e-07 V_hig
+ 3.877010000e-07 V_hig
+ 3.878000000e-07 V_hig
+ 3.878010000e-07 V_hig
+ 3.879000000e-07 V_hig
+ 3.879010000e-07 V_low
+ 3.880000000e-07 V_low
+ 3.880010000e-07 V_low
+ 3.881000000e-07 V_low
+ 3.881010000e-07 V_low
+ 3.882000000e-07 V_low
+ 3.882010000e-07 V_low
+ 3.883000000e-07 V_low
+ 3.883010000e-07 V_low
+ 3.884000000e-07 V_low
+ 3.884010000e-07 V_low
+ 3.885000000e-07 V_low
+ 3.885010000e-07 V_low
+ 3.886000000e-07 V_low
+ 3.886010000e-07 V_low
+ 3.887000000e-07 V_low
+ 3.887010000e-07 V_low
+ 3.888000000e-07 V_low
+ 3.888010000e-07 V_low
+ 3.889000000e-07 V_low
+ 3.889010000e-07 V_low
+ 3.890000000e-07 V_low
+ 3.890010000e-07 V_low
+ 3.891000000e-07 V_low
+ 3.891010000e-07 V_low
+ 3.892000000e-07 V_low
+ 3.892010000e-07 V_low
+ 3.893000000e-07 V_low
+ 3.893010000e-07 V_low
+ 3.894000000e-07 V_low
+ 3.894010000e-07 V_low
+ 3.895000000e-07 V_low
+ 3.895010000e-07 V_low
+ 3.896000000e-07 V_low
+ 3.896010000e-07 V_low
+ 3.897000000e-07 V_low
+ 3.897010000e-07 V_low
+ 3.898000000e-07 V_low
+ 3.898010000e-07 V_low
+ 3.899000000e-07 V_low
+ 3.899010000e-07 V_hig
+ 3.900000000e-07 V_hig
+ 3.900010000e-07 V_hig
+ 3.901000000e-07 V_hig
+ 3.901010000e-07 V_hig
+ 3.902000000e-07 V_hig
+ 3.902010000e-07 V_hig
+ 3.903000000e-07 V_hig
+ 3.903010000e-07 V_hig
+ 3.904000000e-07 V_hig
+ 3.904010000e-07 V_hig
+ 3.905000000e-07 V_hig
+ 3.905010000e-07 V_hig
+ 3.906000000e-07 V_hig
+ 3.906010000e-07 V_hig
+ 3.907000000e-07 V_hig
+ 3.907010000e-07 V_hig
+ 3.908000000e-07 V_hig
+ 3.908010000e-07 V_hig
+ 3.909000000e-07 V_hig
+ 3.909010000e-07 V_low
+ 3.910000000e-07 V_low
+ 3.910010000e-07 V_low
+ 3.911000000e-07 V_low
+ 3.911010000e-07 V_low
+ 3.912000000e-07 V_low
+ 3.912010000e-07 V_low
+ 3.913000000e-07 V_low
+ 3.913010000e-07 V_low
+ 3.914000000e-07 V_low
+ 3.914010000e-07 V_low
+ 3.915000000e-07 V_low
+ 3.915010000e-07 V_low
+ 3.916000000e-07 V_low
+ 3.916010000e-07 V_low
+ 3.917000000e-07 V_low
+ 3.917010000e-07 V_low
+ 3.918000000e-07 V_low
+ 3.918010000e-07 V_low
+ 3.919000000e-07 V_low
+ 3.919010000e-07 V_low
+ 3.920000000e-07 V_low
+ 3.920010000e-07 V_low
+ 3.921000000e-07 V_low
+ 3.921010000e-07 V_low
+ 3.922000000e-07 V_low
+ 3.922010000e-07 V_low
+ 3.923000000e-07 V_low
+ 3.923010000e-07 V_low
+ 3.924000000e-07 V_low
+ 3.924010000e-07 V_low
+ 3.925000000e-07 V_low
+ 3.925010000e-07 V_low
+ 3.926000000e-07 V_low
+ 3.926010000e-07 V_low
+ 3.927000000e-07 V_low
+ 3.927010000e-07 V_low
+ 3.928000000e-07 V_low
+ 3.928010000e-07 V_low
+ 3.929000000e-07 V_low
+ 3.929010000e-07 V_hig
+ 3.930000000e-07 V_hig
+ 3.930010000e-07 V_hig
+ 3.931000000e-07 V_hig
+ 3.931010000e-07 V_hig
+ 3.932000000e-07 V_hig
+ 3.932010000e-07 V_hig
+ 3.933000000e-07 V_hig
+ 3.933010000e-07 V_hig
+ 3.934000000e-07 V_hig
+ 3.934010000e-07 V_hig
+ 3.935000000e-07 V_hig
+ 3.935010000e-07 V_hig
+ 3.936000000e-07 V_hig
+ 3.936010000e-07 V_hig
+ 3.937000000e-07 V_hig
+ 3.937010000e-07 V_hig
+ 3.938000000e-07 V_hig
+ 3.938010000e-07 V_hig
+ 3.939000000e-07 V_hig
+ 3.939010000e-07 V_low
+ 3.940000000e-07 V_low
+ 3.940010000e-07 V_low
+ 3.941000000e-07 V_low
+ 3.941010000e-07 V_low
+ 3.942000000e-07 V_low
+ 3.942010000e-07 V_low
+ 3.943000000e-07 V_low
+ 3.943010000e-07 V_low
+ 3.944000000e-07 V_low
+ 3.944010000e-07 V_low
+ 3.945000000e-07 V_low
+ 3.945010000e-07 V_low
+ 3.946000000e-07 V_low
+ 3.946010000e-07 V_low
+ 3.947000000e-07 V_low
+ 3.947010000e-07 V_low
+ 3.948000000e-07 V_low
+ 3.948010000e-07 V_low
+ 3.949000000e-07 V_low
+ 3.949010000e-07 V_hig
+ 3.950000000e-07 V_hig
+ 3.950010000e-07 V_hig
+ 3.951000000e-07 V_hig
+ 3.951010000e-07 V_hig
+ 3.952000000e-07 V_hig
+ 3.952010000e-07 V_hig
+ 3.953000000e-07 V_hig
+ 3.953010000e-07 V_hig
+ 3.954000000e-07 V_hig
+ 3.954010000e-07 V_hig
+ 3.955000000e-07 V_hig
+ 3.955010000e-07 V_hig
+ 3.956000000e-07 V_hig
+ 3.956010000e-07 V_hig
+ 3.957000000e-07 V_hig
+ 3.957010000e-07 V_hig
+ 3.958000000e-07 V_hig
+ 3.958010000e-07 V_hig
+ 3.959000000e-07 V_hig
+ 3.959010000e-07 V_hig
+ 3.960000000e-07 V_hig
+ 3.960010000e-07 V_hig
+ 3.961000000e-07 V_hig
+ 3.961010000e-07 V_hig
+ 3.962000000e-07 V_hig
+ 3.962010000e-07 V_hig
+ 3.963000000e-07 V_hig
+ 3.963010000e-07 V_hig
+ 3.964000000e-07 V_hig
+ 3.964010000e-07 V_hig
+ 3.965000000e-07 V_hig
+ 3.965010000e-07 V_hig
+ 3.966000000e-07 V_hig
+ 3.966010000e-07 V_hig
+ 3.967000000e-07 V_hig
+ 3.967010000e-07 V_hig
+ 3.968000000e-07 V_hig
+ 3.968010000e-07 V_hig
+ 3.969000000e-07 V_hig
+ 3.969010000e-07 V_low
+ 3.970000000e-07 V_low
+ 3.970010000e-07 V_low
+ 3.971000000e-07 V_low
+ 3.971010000e-07 V_low
+ 3.972000000e-07 V_low
+ 3.972010000e-07 V_low
+ 3.973000000e-07 V_low
+ 3.973010000e-07 V_low
+ 3.974000000e-07 V_low
+ 3.974010000e-07 V_low
+ 3.975000000e-07 V_low
+ 3.975010000e-07 V_low
+ 3.976000000e-07 V_low
+ 3.976010000e-07 V_low
+ 3.977000000e-07 V_low
+ 3.977010000e-07 V_low
+ 3.978000000e-07 V_low
+ 3.978010000e-07 V_low
+ 3.979000000e-07 V_low
+ 3.979010000e-07 V_hig
+ 3.980000000e-07 V_hig
+ 3.980010000e-07 V_hig
+ 3.981000000e-07 V_hig
+ 3.981010000e-07 V_hig
+ 3.982000000e-07 V_hig
+ 3.982010000e-07 V_hig
+ 3.983000000e-07 V_hig
+ 3.983010000e-07 V_hig
+ 3.984000000e-07 V_hig
+ 3.984010000e-07 V_hig
+ 3.985000000e-07 V_hig
+ 3.985010000e-07 V_hig
+ 3.986000000e-07 V_hig
+ 3.986010000e-07 V_hig
+ 3.987000000e-07 V_hig
+ 3.987010000e-07 V_hig
+ 3.988000000e-07 V_hig
+ 3.988010000e-07 V_hig
+ 3.989000000e-07 V_hig
+ 3.989010000e-07 V_hig
+ 3.990000000e-07 V_hig
+ 3.990010000e-07 V_hig
+ 3.991000000e-07 V_hig
+ 3.991010000e-07 V_hig
+ 3.992000000e-07 V_hig
+ 3.992010000e-07 V_hig
+ 3.993000000e-07 V_hig
+ 3.993010000e-07 V_hig
+ 3.994000000e-07 V_hig
+ 3.994010000e-07 V_hig
+ 3.995000000e-07 V_hig
+ 3.995010000e-07 V_hig
+ 3.996000000e-07 V_hig
+ 3.996010000e-07 V_hig
+ 3.997000000e-07 V_hig
+ 3.997010000e-07 V_hig
+ 3.998000000e-07 V_hig
+ 3.998010000e-07 V_hig
+ 3.999000000e-07 V_hig
+ 3.999010000e-07 V_hig
+ 4.000000000e-07 V_hig
+ 4.000010000e-07 V_hig
+ 4.001000000e-07 V_hig
+ 4.001010000e-07 V_hig
+ 4.002000000e-07 V_hig
+ 4.002010000e-07 V_hig
+ 4.003000000e-07 V_hig
+ 4.003010000e-07 V_hig
+ 4.004000000e-07 V_hig
+ 4.004010000e-07 V_hig
+ 4.005000000e-07 V_hig
+ 4.005010000e-07 V_hig
+ 4.006000000e-07 V_hig
+ 4.006010000e-07 V_hig
+ 4.007000000e-07 V_hig
+ 4.007010000e-07 V_hig
+ 4.008000000e-07 V_hig
+ 4.008010000e-07 V_hig
+ 4.009000000e-07 V_hig
+ 4.009010000e-07 V_low
+ 4.010000000e-07 V_low
+ 4.010010000e-07 V_low
+ 4.011000000e-07 V_low
+ 4.011010000e-07 V_low
+ 4.012000000e-07 V_low
+ 4.012010000e-07 V_low
+ 4.013000000e-07 V_low
+ 4.013010000e-07 V_low
+ 4.014000000e-07 V_low
+ 4.014010000e-07 V_low
+ 4.015000000e-07 V_low
+ 4.015010000e-07 V_low
+ 4.016000000e-07 V_low
+ 4.016010000e-07 V_low
+ 4.017000000e-07 V_low
+ 4.017010000e-07 V_low
+ 4.018000000e-07 V_low
+ 4.018010000e-07 V_low
+ 4.019000000e-07 V_low
+ 4.019010000e-07 V_hig
+ 4.020000000e-07 V_hig
+ 4.020010000e-07 V_hig
+ 4.021000000e-07 V_hig
+ 4.021010000e-07 V_hig
+ 4.022000000e-07 V_hig
+ 4.022010000e-07 V_hig
+ 4.023000000e-07 V_hig
+ 4.023010000e-07 V_hig
+ 4.024000000e-07 V_hig
+ 4.024010000e-07 V_hig
+ 4.025000000e-07 V_hig
+ 4.025010000e-07 V_hig
+ 4.026000000e-07 V_hig
+ 4.026010000e-07 V_hig
+ 4.027000000e-07 V_hig
+ 4.027010000e-07 V_hig
+ 4.028000000e-07 V_hig
+ 4.028010000e-07 V_hig
+ 4.029000000e-07 V_hig
+ 4.029010000e-07 V_hig
+ 4.030000000e-07 V_hig
+ 4.030010000e-07 V_hig
+ 4.031000000e-07 V_hig
+ 4.031010000e-07 V_hig
+ 4.032000000e-07 V_hig
+ 4.032010000e-07 V_hig
+ 4.033000000e-07 V_hig
+ 4.033010000e-07 V_hig
+ 4.034000000e-07 V_hig
+ 4.034010000e-07 V_hig
+ 4.035000000e-07 V_hig
+ 4.035010000e-07 V_hig
+ 4.036000000e-07 V_hig
+ 4.036010000e-07 V_hig
+ 4.037000000e-07 V_hig
+ 4.037010000e-07 V_hig
+ 4.038000000e-07 V_hig
+ 4.038010000e-07 V_hig
+ 4.039000000e-07 V_hig
+ 4.039010000e-07 V_low
+ 4.040000000e-07 V_low
+ 4.040010000e-07 V_low
+ 4.041000000e-07 V_low
+ 4.041010000e-07 V_low
+ 4.042000000e-07 V_low
+ 4.042010000e-07 V_low
+ 4.043000000e-07 V_low
+ 4.043010000e-07 V_low
+ 4.044000000e-07 V_low
+ 4.044010000e-07 V_low
+ 4.045000000e-07 V_low
+ 4.045010000e-07 V_low
+ 4.046000000e-07 V_low
+ 4.046010000e-07 V_low
+ 4.047000000e-07 V_low
+ 4.047010000e-07 V_low
+ 4.048000000e-07 V_low
+ 4.048010000e-07 V_low
+ 4.049000000e-07 V_low
+ 4.049010000e-07 V_low
+ 4.050000000e-07 V_low
+ 4.050010000e-07 V_low
+ 4.051000000e-07 V_low
+ 4.051010000e-07 V_low
+ 4.052000000e-07 V_low
+ 4.052010000e-07 V_low
+ 4.053000000e-07 V_low
+ 4.053010000e-07 V_low
+ 4.054000000e-07 V_low
+ 4.054010000e-07 V_low
+ 4.055000000e-07 V_low
+ 4.055010000e-07 V_low
+ 4.056000000e-07 V_low
+ 4.056010000e-07 V_low
+ 4.057000000e-07 V_low
+ 4.057010000e-07 V_low
+ 4.058000000e-07 V_low
+ 4.058010000e-07 V_low
+ 4.059000000e-07 V_low
+ 4.059010000e-07 V_low
+ 4.060000000e-07 V_low
+ 4.060010000e-07 V_low
+ 4.061000000e-07 V_low
+ 4.061010000e-07 V_low
+ 4.062000000e-07 V_low
+ 4.062010000e-07 V_low
+ 4.063000000e-07 V_low
+ 4.063010000e-07 V_low
+ 4.064000000e-07 V_low
+ 4.064010000e-07 V_low
+ 4.065000000e-07 V_low
+ 4.065010000e-07 V_low
+ 4.066000000e-07 V_low
+ 4.066010000e-07 V_low
+ 4.067000000e-07 V_low
+ 4.067010000e-07 V_low
+ 4.068000000e-07 V_low
+ 4.068010000e-07 V_low
+ 4.069000000e-07 V_low
+ 4.069010000e-07 V_low
+ 4.070000000e-07 V_low
+ 4.070010000e-07 V_low
+ 4.071000000e-07 V_low
+ 4.071010000e-07 V_low
+ 4.072000000e-07 V_low
+ 4.072010000e-07 V_low
+ 4.073000000e-07 V_low
+ 4.073010000e-07 V_low
+ 4.074000000e-07 V_low
+ 4.074010000e-07 V_low
+ 4.075000000e-07 V_low
+ 4.075010000e-07 V_low
+ 4.076000000e-07 V_low
+ 4.076010000e-07 V_low
+ 4.077000000e-07 V_low
+ 4.077010000e-07 V_low
+ 4.078000000e-07 V_low
+ 4.078010000e-07 V_low
+ 4.079000000e-07 V_low
+ 4.079010000e-07 V_hig
+ 4.080000000e-07 V_hig
+ 4.080010000e-07 V_hig
+ 4.081000000e-07 V_hig
+ 4.081010000e-07 V_hig
+ 4.082000000e-07 V_hig
+ 4.082010000e-07 V_hig
+ 4.083000000e-07 V_hig
+ 4.083010000e-07 V_hig
+ 4.084000000e-07 V_hig
+ 4.084010000e-07 V_hig
+ 4.085000000e-07 V_hig
+ 4.085010000e-07 V_hig
+ 4.086000000e-07 V_hig
+ 4.086010000e-07 V_hig
+ 4.087000000e-07 V_hig
+ 4.087010000e-07 V_hig
+ 4.088000000e-07 V_hig
+ 4.088010000e-07 V_hig
+ 4.089000000e-07 V_hig
+ 4.089010000e-07 V_hig
+ 4.090000000e-07 V_hig
+ 4.090010000e-07 V_hig
+ 4.091000000e-07 V_hig
+ 4.091010000e-07 V_hig
+ 4.092000000e-07 V_hig
+ 4.092010000e-07 V_hig
+ 4.093000000e-07 V_hig
+ 4.093010000e-07 V_hig
+ 4.094000000e-07 V_hig
+ 4.094010000e-07 V_hig
+ 4.095000000e-07 V_hig
+ 4.095010000e-07 V_hig
+ 4.096000000e-07 V_hig
+ 4.096010000e-07 V_hig
+ 4.097000000e-07 V_hig
+ 4.097010000e-07 V_hig
+ 4.098000000e-07 V_hig
+ 4.098010000e-07 V_hig
+ 4.099000000e-07 V_hig
+ 4.099010000e-07 V_hig
+ 4.100000000e-07 V_hig
+ 4.100010000e-07 V_hig
+ 4.101000000e-07 V_hig
+ 4.101010000e-07 V_hig
+ 4.102000000e-07 V_hig
+ 4.102010000e-07 V_hig
+ 4.103000000e-07 V_hig
+ 4.103010000e-07 V_hig
+ 4.104000000e-07 V_hig
+ 4.104010000e-07 V_hig
+ 4.105000000e-07 V_hig
+ 4.105010000e-07 V_hig
+ 4.106000000e-07 V_hig
+ 4.106010000e-07 V_hig
+ 4.107000000e-07 V_hig
+ 4.107010000e-07 V_hig
+ 4.108000000e-07 V_hig
+ 4.108010000e-07 V_hig
+ 4.109000000e-07 V_hig
+ 4.109010000e-07 V_hig
+ 4.110000000e-07 V_hig
+ 4.110010000e-07 V_hig
+ 4.111000000e-07 V_hig
+ 4.111010000e-07 V_hig
+ 4.112000000e-07 V_hig
+ 4.112010000e-07 V_hig
+ 4.113000000e-07 V_hig
+ 4.113010000e-07 V_hig
+ 4.114000000e-07 V_hig
+ 4.114010000e-07 V_hig
+ 4.115000000e-07 V_hig
+ 4.115010000e-07 V_hig
+ 4.116000000e-07 V_hig
+ 4.116010000e-07 V_hig
+ 4.117000000e-07 V_hig
+ 4.117010000e-07 V_hig
+ 4.118000000e-07 V_hig
+ 4.118010000e-07 V_hig
+ 4.119000000e-07 V_hig
+ 4.119010000e-07 V_low
+ 4.120000000e-07 V_low
+ 4.120010000e-07 V_low
+ 4.121000000e-07 V_low
+ 4.121010000e-07 V_low
+ 4.122000000e-07 V_low
+ 4.122010000e-07 V_low
+ 4.123000000e-07 V_low
+ 4.123010000e-07 V_low
+ 4.124000000e-07 V_low
+ 4.124010000e-07 V_low
+ 4.125000000e-07 V_low
+ 4.125010000e-07 V_low
+ 4.126000000e-07 V_low
+ 4.126010000e-07 V_low
+ 4.127000000e-07 V_low
+ 4.127010000e-07 V_low
+ 4.128000000e-07 V_low
+ 4.128010000e-07 V_low
+ 4.129000000e-07 V_low
+ 4.129010000e-07 V_low
+ 4.130000000e-07 V_low
+ 4.130010000e-07 V_low
+ 4.131000000e-07 V_low
+ 4.131010000e-07 V_low
+ 4.132000000e-07 V_low
+ 4.132010000e-07 V_low
+ 4.133000000e-07 V_low
+ 4.133010000e-07 V_low
+ 4.134000000e-07 V_low
+ 4.134010000e-07 V_low
+ 4.135000000e-07 V_low
+ 4.135010000e-07 V_low
+ 4.136000000e-07 V_low
+ 4.136010000e-07 V_low
+ 4.137000000e-07 V_low
+ 4.137010000e-07 V_low
+ 4.138000000e-07 V_low
+ 4.138010000e-07 V_low
+ 4.139000000e-07 V_low
+ 4.139010000e-07 V_hig
+ 4.140000000e-07 V_hig
+ 4.140010000e-07 V_hig
+ 4.141000000e-07 V_hig
+ 4.141010000e-07 V_hig
+ 4.142000000e-07 V_hig
+ 4.142010000e-07 V_hig
+ 4.143000000e-07 V_hig
+ 4.143010000e-07 V_hig
+ 4.144000000e-07 V_hig
+ 4.144010000e-07 V_hig
+ 4.145000000e-07 V_hig
+ 4.145010000e-07 V_hig
+ 4.146000000e-07 V_hig
+ 4.146010000e-07 V_hig
+ 4.147000000e-07 V_hig
+ 4.147010000e-07 V_hig
+ 4.148000000e-07 V_hig
+ 4.148010000e-07 V_hig
+ 4.149000000e-07 V_hig
+ 4.149010000e-07 V_hig
+ 4.150000000e-07 V_hig
+ 4.150010000e-07 V_hig
+ 4.151000000e-07 V_hig
+ 4.151010000e-07 V_hig
+ 4.152000000e-07 V_hig
+ 4.152010000e-07 V_hig
+ 4.153000000e-07 V_hig
+ 4.153010000e-07 V_hig
+ 4.154000000e-07 V_hig
+ 4.154010000e-07 V_hig
+ 4.155000000e-07 V_hig
+ 4.155010000e-07 V_hig
+ 4.156000000e-07 V_hig
+ 4.156010000e-07 V_hig
+ 4.157000000e-07 V_hig
+ 4.157010000e-07 V_hig
+ 4.158000000e-07 V_hig
+ 4.158010000e-07 V_hig
+ 4.159000000e-07 V_hig
+ 4.159010000e-07 V_low
+ 4.160000000e-07 V_low
+ 4.160010000e-07 V_low
+ 4.161000000e-07 V_low
+ 4.161010000e-07 V_low
+ 4.162000000e-07 V_low
+ 4.162010000e-07 V_low
+ 4.163000000e-07 V_low
+ 4.163010000e-07 V_low
+ 4.164000000e-07 V_low
+ 4.164010000e-07 V_low
+ 4.165000000e-07 V_low
+ 4.165010000e-07 V_low
+ 4.166000000e-07 V_low
+ 4.166010000e-07 V_low
+ 4.167000000e-07 V_low
+ 4.167010000e-07 V_low
+ 4.168000000e-07 V_low
+ 4.168010000e-07 V_low
+ 4.169000000e-07 V_low
+ 4.169010000e-07 V_hig
+ 4.170000000e-07 V_hig
+ 4.170010000e-07 V_hig
+ 4.171000000e-07 V_hig
+ 4.171010000e-07 V_hig
+ 4.172000000e-07 V_hig
+ 4.172010000e-07 V_hig
+ 4.173000000e-07 V_hig
+ 4.173010000e-07 V_hig
+ 4.174000000e-07 V_hig
+ 4.174010000e-07 V_hig
+ 4.175000000e-07 V_hig
+ 4.175010000e-07 V_hig
+ 4.176000000e-07 V_hig
+ 4.176010000e-07 V_hig
+ 4.177000000e-07 V_hig
+ 4.177010000e-07 V_hig
+ 4.178000000e-07 V_hig
+ 4.178010000e-07 V_hig
+ 4.179000000e-07 V_hig
+ 4.179010000e-07 V_hig
+ 4.180000000e-07 V_hig
+ 4.180010000e-07 V_hig
+ 4.181000000e-07 V_hig
+ 4.181010000e-07 V_hig
+ 4.182000000e-07 V_hig
+ 4.182010000e-07 V_hig
+ 4.183000000e-07 V_hig
+ 4.183010000e-07 V_hig
+ 4.184000000e-07 V_hig
+ 4.184010000e-07 V_hig
+ 4.185000000e-07 V_hig
+ 4.185010000e-07 V_hig
+ 4.186000000e-07 V_hig
+ 4.186010000e-07 V_hig
+ 4.187000000e-07 V_hig
+ 4.187010000e-07 V_hig
+ 4.188000000e-07 V_hig
+ 4.188010000e-07 V_hig
+ 4.189000000e-07 V_hig
+ 4.189010000e-07 V_low
+ 4.190000000e-07 V_low
+ 4.190010000e-07 V_low
+ 4.191000000e-07 V_low
+ 4.191010000e-07 V_low
+ 4.192000000e-07 V_low
+ 4.192010000e-07 V_low
+ 4.193000000e-07 V_low
+ 4.193010000e-07 V_low
+ 4.194000000e-07 V_low
+ 4.194010000e-07 V_low
+ 4.195000000e-07 V_low
+ 4.195010000e-07 V_low
+ 4.196000000e-07 V_low
+ 4.196010000e-07 V_low
+ 4.197000000e-07 V_low
+ 4.197010000e-07 V_low
+ 4.198000000e-07 V_low
+ 4.198010000e-07 V_low
+ 4.199000000e-07 V_low
+ 4.199010000e-07 V_hig
+ 4.200000000e-07 V_hig
+ 4.200010000e-07 V_hig
+ 4.201000000e-07 V_hig
+ 4.201010000e-07 V_hig
+ 4.202000000e-07 V_hig
+ 4.202010000e-07 V_hig
+ 4.203000000e-07 V_hig
+ 4.203010000e-07 V_hig
+ 4.204000000e-07 V_hig
+ 4.204010000e-07 V_hig
+ 4.205000000e-07 V_hig
+ 4.205010000e-07 V_hig
+ 4.206000000e-07 V_hig
+ 4.206010000e-07 V_hig
+ 4.207000000e-07 V_hig
+ 4.207010000e-07 V_hig
+ 4.208000000e-07 V_hig
+ 4.208010000e-07 V_hig
+ 4.209000000e-07 V_hig
+ 4.209010000e-07 V_hig
+ 4.210000000e-07 V_hig
+ 4.210010000e-07 V_hig
+ 4.211000000e-07 V_hig
+ 4.211010000e-07 V_hig
+ 4.212000000e-07 V_hig
+ 4.212010000e-07 V_hig
+ 4.213000000e-07 V_hig
+ 4.213010000e-07 V_hig
+ 4.214000000e-07 V_hig
+ 4.214010000e-07 V_hig
+ 4.215000000e-07 V_hig
+ 4.215010000e-07 V_hig
+ 4.216000000e-07 V_hig
+ 4.216010000e-07 V_hig
+ 4.217000000e-07 V_hig
+ 4.217010000e-07 V_hig
+ 4.218000000e-07 V_hig
+ 4.218010000e-07 V_hig
+ 4.219000000e-07 V_hig
+ 4.219010000e-07 V_hig
+ 4.220000000e-07 V_hig
+ 4.220010000e-07 V_hig
+ 4.221000000e-07 V_hig
+ 4.221010000e-07 V_hig
+ 4.222000000e-07 V_hig
+ 4.222010000e-07 V_hig
+ 4.223000000e-07 V_hig
+ 4.223010000e-07 V_hig
+ 4.224000000e-07 V_hig
+ 4.224010000e-07 V_hig
+ 4.225000000e-07 V_hig
+ 4.225010000e-07 V_hig
+ 4.226000000e-07 V_hig
+ 4.226010000e-07 V_hig
+ 4.227000000e-07 V_hig
+ 4.227010000e-07 V_hig
+ 4.228000000e-07 V_hig
+ 4.228010000e-07 V_hig
+ 4.229000000e-07 V_hig
+ 4.229010000e-07 V_hig
+ 4.230000000e-07 V_hig
+ 4.230010000e-07 V_hig
+ 4.231000000e-07 V_hig
+ 4.231010000e-07 V_hig
+ 4.232000000e-07 V_hig
+ 4.232010000e-07 V_hig
+ 4.233000000e-07 V_hig
+ 4.233010000e-07 V_hig
+ 4.234000000e-07 V_hig
+ 4.234010000e-07 V_hig
+ 4.235000000e-07 V_hig
+ 4.235010000e-07 V_hig
+ 4.236000000e-07 V_hig
+ 4.236010000e-07 V_hig
+ 4.237000000e-07 V_hig
+ 4.237010000e-07 V_hig
+ 4.238000000e-07 V_hig
+ 4.238010000e-07 V_hig
+ 4.239000000e-07 V_hig
+ 4.239010000e-07 V_hig
+ 4.240000000e-07 V_hig
+ 4.240010000e-07 V_hig
+ 4.241000000e-07 V_hig
+ 4.241010000e-07 V_hig
+ 4.242000000e-07 V_hig
+ 4.242010000e-07 V_hig
+ 4.243000000e-07 V_hig
+ 4.243010000e-07 V_hig
+ 4.244000000e-07 V_hig
+ 4.244010000e-07 V_hig
+ 4.245000000e-07 V_hig
+ 4.245010000e-07 V_hig
+ 4.246000000e-07 V_hig
+ 4.246010000e-07 V_hig
+ 4.247000000e-07 V_hig
+ 4.247010000e-07 V_hig
+ 4.248000000e-07 V_hig
+ 4.248010000e-07 V_hig
+ 4.249000000e-07 V_hig
+ 4.249010000e-07 V_hig
+ 4.250000000e-07 V_hig
+ 4.250010000e-07 V_hig
+ 4.251000000e-07 V_hig
+ 4.251010000e-07 V_hig
+ 4.252000000e-07 V_hig
+ 4.252010000e-07 V_hig
+ 4.253000000e-07 V_hig
+ 4.253010000e-07 V_hig
+ 4.254000000e-07 V_hig
+ 4.254010000e-07 V_hig
+ 4.255000000e-07 V_hig
+ 4.255010000e-07 V_hig
+ 4.256000000e-07 V_hig
+ 4.256010000e-07 V_hig
+ 4.257000000e-07 V_hig
+ 4.257010000e-07 V_hig
+ 4.258000000e-07 V_hig
+ 4.258010000e-07 V_hig
+ 4.259000000e-07 V_hig
+ 4.259010000e-07 V_hig
+ 4.260000000e-07 V_hig
+ 4.260010000e-07 V_hig
+ 4.261000000e-07 V_hig
+ 4.261010000e-07 V_hig
+ 4.262000000e-07 V_hig
+ 4.262010000e-07 V_hig
+ 4.263000000e-07 V_hig
+ 4.263010000e-07 V_hig
+ 4.264000000e-07 V_hig
+ 4.264010000e-07 V_hig
+ 4.265000000e-07 V_hig
+ 4.265010000e-07 V_hig
+ 4.266000000e-07 V_hig
+ 4.266010000e-07 V_hig
+ 4.267000000e-07 V_hig
+ 4.267010000e-07 V_hig
+ 4.268000000e-07 V_hig
+ 4.268010000e-07 V_hig
+ 4.269000000e-07 V_hig
+ 4.269010000e-07 V_low
+ 4.270000000e-07 V_low
+ 4.270010000e-07 V_low
+ 4.271000000e-07 V_low
+ 4.271010000e-07 V_low
+ 4.272000000e-07 V_low
+ 4.272010000e-07 V_low
+ 4.273000000e-07 V_low
+ 4.273010000e-07 V_low
+ 4.274000000e-07 V_low
+ 4.274010000e-07 V_low
+ 4.275000000e-07 V_low
+ 4.275010000e-07 V_low
+ 4.276000000e-07 V_low
+ 4.276010000e-07 V_low
+ 4.277000000e-07 V_low
+ 4.277010000e-07 V_low
+ 4.278000000e-07 V_low
+ 4.278010000e-07 V_low
+ 4.279000000e-07 V_low
+ 4.279010000e-07 V_hig
+ 4.280000000e-07 V_hig
+ 4.280010000e-07 V_hig
+ 4.281000000e-07 V_hig
+ 4.281010000e-07 V_hig
+ 4.282000000e-07 V_hig
+ 4.282010000e-07 V_hig
+ 4.283000000e-07 V_hig
+ 4.283010000e-07 V_hig
+ 4.284000000e-07 V_hig
+ 4.284010000e-07 V_hig
+ 4.285000000e-07 V_hig
+ 4.285010000e-07 V_hig
+ 4.286000000e-07 V_hig
+ 4.286010000e-07 V_hig
+ 4.287000000e-07 V_hig
+ 4.287010000e-07 V_hig
+ 4.288000000e-07 V_hig
+ 4.288010000e-07 V_hig
+ 4.289000000e-07 V_hig
+ 4.289010000e-07 V_hig
+ 4.290000000e-07 V_hig
+ 4.290010000e-07 V_hig
+ 4.291000000e-07 V_hig
+ 4.291010000e-07 V_hig
+ 4.292000000e-07 V_hig
+ 4.292010000e-07 V_hig
+ 4.293000000e-07 V_hig
+ 4.293010000e-07 V_hig
+ 4.294000000e-07 V_hig
+ 4.294010000e-07 V_hig
+ 4.295000000e-07 V_hig
+ 4.295010000e-07 V_hig
+ 4.296000000e-07 V_hig
+ 4.296010000e-07 V_hig
+ 4.297000000e-07 V_hig
+ 4.297010000e-07 V_hig
+ 4.298000000e-07 V_hig
+ 4.298010000e-07 V_hig
+ 4.299000000e-07 V_hig
+ 4.299010000e-07 V_hig
+ 4.300000000e-07 V_hig
+ 4.300010000e-07 V_hig
+ 4.301000000e-07 V_hig
+ 4.301010000e-07 V_hig
+ 4.302000000e-07 V_hig
+ 4.302010000e-07 V_hig
+ 4.303000000e-07 V_hig
+ 4.303010000e-07 V_hig
+ 4.304000000e-07 V_hig
+ 4.304010000e-07 V_hig
+ 4.305000000e-07 V_hig
+ 4.305010000e-07 V_hig
+ 4.306000000e-07 V_hig
+ 4.306010000e-07 V_hig
+ 4.307000000e-07 V_hig
+ 4.307010000e-07 V_hig
+ 4.308000000e-07 V_hig
+ 4.308010000e-07 V_hig
+ 4.309000000e-07 V_hig
+ 4.309010000e-07 V_low
+ 4.310000000e-07 V_low
+ 4.310010000e-07 V_low
+ 4.311000000e-07 V_low
+ 4.311010000e-07 V_low
+ 4.312000000e-07 V_low
+ 4.312010000e-07 V_low
+ 4.313000000e-07 V_low
+ 4.313010000e-07 V_low
+ 4.314000000e-07 V_low
+ 4.314010000e-07 V_low
+ 4.315000000e-07 V_low
+ 4.315010000e-07 V_low
+ 4.316000000e-07 V_low
+ 4.316010000e-07 V_low
+ 4.317000000e-07 V_low
+ 4.317010000e-07 V_low
+ 4.318000000e-07 V_low
+ 4.318010000e-07 V_low
+ 4.319000000e-07 V_low
+ 4.319010000e-07 V_low
+ 4.320000000e-07 V_low
+ 4.320010000e-07 V_low
+ 4.321000000e-07 V_low
+ 4.321010000e-07 V_low
+ 4.322000000e-07 V_low
+ 4.322010000e-07 V_low
+ 4.323000000e-07 V_low
+ 4.323010000e-07 V_low
+ 4.324000000e-07 V_low
+ 4.324010000e-07 V_low
+ 4.325000000e-07 V_low
+ 4.325010000e-07 V_low
+ 4.326000000e-07 V_low
+ 4.326010000e-07 V_low
+ 4.327000000e-07 V_low
+ 4.327010000e-07 V_low
+ 4.328000000e-07 V_low
+ 4.328010000e-07 V_low
+ 4.329000000e-07 V_low
+ 4.329010000e-07 V_low
+ 4.330000000e-07 V_low
+ 4.330010000e-07 V_low
+ 4.331000000e-07 V_low
+ 4.331010000e-07 V_low
+ 4.332000000e-07 V_low
+ 4.332010000e-07 V_low
+ 4.333000000e-07 V_low
+ 4.333010000e-07 V_low
+ 4.334000000e-07 V_low
+ 4.334010000e-07 V_low
+ 4.335000000e-07 V_low
+ 4.335010000e-07 V_low
+ 4.336000000e-07 V_low
+ 4.336010000e-07 V_low
+ 4.337000000e-07 V_low
+ 4.337010000e-07 V_low
+ 4.338000000e-07 V_low
+ 4.338010000e-07 V_low
+ 4.339000000e-07 V_low
+ 4.339010000e-07 V_hig
+ 4.340000000e-07 V_hig
+ 4.340010000e-07 V_hig
+ 4.341000000e-07 V_hig
+ 4.341010000e-07 V_hig
+ 4.342000000e-07 V_hig
+ 4.342010000e-07 V_hig
+ 4.343000000e-07 V_hig
+ 4.343010000e-07 V_hig
+ 4.344000000e-07 V_hig
+ 4.344010000e-07 V_hig
+ 4.345000000e-07 V_hig
+ 4.345010000e-07 V_hig
+ 4.346000000e-07 V_hig
+ 4.346010000e-07 V_hig
+ 4.347000000e-07 V_hig
+ 4.347010000e-07 V_hig
+ 4.348000000e-07 V_hig
+ 4.348010000e-07 V_hig
+ 4.349000000e-07 V_hig
+ 4.349010000e-07 V_low
+ 4.350000000e-07 V_low
+ 4.350010000e-07 V_low
+ 4.351000000e-07 V_low
+ 4.351010000e-07 V_low
+ 4.352000000e-07 V_low
+ 4.352010000e-07 V_low
+ 4.353000000e-07 V_low
+ 4.353010000e-07 V_low
+ 4.354000000e-07 V_low
+ 4.354010000e-07 V_low
+ 4.355000000e-07 V_low
+ 4.355010000e-07 V_low
+ 4.356000000e-07 V_low
+ 4.356010000e-07 V_low
+ 4.357000000e-07 V_low
+ 4.357010000e-07 V_low
+ 4.358000000e-07 V_low
+ 4.358010000e-07 V_low
+ 4.359000000e-07 V_low
+ 4.359010000e-07 V_hig
+ 4.360000000e-07 V_hig
+ 4.360010000e-07 V_hig
+ 4.361000000e-07 V_hig
+ 4.361010000e-07 V_hig
+ 4.362000000e-07 V_hig
+ 4.362010000e-07 V_hig
+ 4.363000000e-07 V_hig
+ 4.363010000e-07 V_hig
+ 4.364000000e-07 V_hig
+ 4.364010000e-07 V_hig
+ 4.365000000e-07 V_hig
+ 4.365010000e-07 V_hig
+ 4.366000000e-07 V_hig
+ 4.366010000e-07 V_hig
+ 4.367000000e-07 V_hig
+ 4.367010000e-07 V_hig
+ 4.368000000e-07 V_hig
+ 4.368010000e-07 V_hig
+ 4.369000000e-07 V_hig
+ 4.369010000e-07 V_hig
+ 4.370000000e-07 V_hig
+ 4.370010000e-07 V_hig
+ 4.371000000e-07 V_hig
+ 4.371010000e-07 V_hig
+ 4.372000000e-07 V_hig
+ 4.372010000e-07 V_hig
+ 4.373000000e-07 V_hig
+ 4.373010000e-07 V_hig
+ 4.374000000e-07 V_hig
+ 4.374010000e-07 V_hig
+ 4.375000000e-07 V_hig
+ 4.375010000e-07 V_hig
+ 4.376000000e-07 V_hig
+ 4.376010000e-07 V_hig
+ 4.377000000e-07 V_hig
+ 4.377010000e-07 V_hig
+ 4.378000000e-07 V_hig
+ 4.378010000e-07 V_hig
+ 4.379000000e-07 V_hig
+ 4.379010000e-07 V_hig
+ 4.380000000e-07 V_hig
+ 4.380010000e-07 V_hig
+ 4.381000000e-07 V_hig
+ 4.381010000e-07 V_hig
+ 4.382000000e-07 V_hig
+ 4.382010000e-07 V_hig
+ 4.383000000e-07 V_hig
+ 4.383010000e-07 V_hig
+ 4.384000000e-07 V_hig
+ 4.384010000e-07 V_hig
+ 4.385000000e-07 V_hig
+ 4.385010000e-07 V_hig
+ 4.386000000e-07 V_hig
+ 4.386010000e-07 V_hig
+ 4.387000000e-07 V_hig
+ 4.387010000e-07 V_hig
+ 4.388000000e-07 V_hig
+ 4.388010000e-07 V_hig
+ 4.389000000e-07 V_hig
+ 4.389010000e-07 V_low
+ 4.390000000e-07 V_low
+ 4.390010000e-07 V_low
+ 4.391000000e-07 V_low
+ 4.391010000e-07 V_low
+ 4.392000000e-07 V_low
+ 4.392010000e-07 V_low
+ 4.393000000e-07 V_low
+ 4.393010000e-07 V_low
+ 4.394000000e-07 V_low
+ 4.394010000e-07 V_low
+ 4.395000000e-07 V_low
+ 4.395010000e-07 V_low
+ 4.396000000e-07 V_low
+ 4.396010000e-07 V_low
+ 4.397000000e-07 V_low
+ 4.397010000e-07 V_low
+ 4.398000000e-07 V_low
+ 4.398010000e-07 V_low
+ 4.399000000e-07 V_low
+ 4.399010000e-07 V_low
+ 4.400000000e-07 V_low
+ 4.400010000e-07 V_low
+ 4.401000000e-07 V_low
+ 4.401010000e-07 V_low
+ 4.402000000e-07 V_low
+ 4.402010000e-07 V_low
+ 4.403000000e-07 V_low
+ 4.403010000e-07 V_low
+ 4.404000000e-07 V_low
+ 4.404010000e-07 V_low
+ 4.405000000e-07 V_low
+ 4.405010000e-07 V_low
+ 4.406000000e-07 V_low
+ 4.406010000e-07 V_low
+ 4.407000000e-07 V_low
+ 4.407010000e-07 V_low
+ 4.408000000e-07 V_low
+ 4.408010000e-07 V_low
+ 4.409000000e-07 V_low
+ 4.409010000e-07 V_low
+ 4.410000000e-07 V_low
+ 4.410010000e-07 V_low
+ 4.411000000e-07 V_low
+ 4.411010000e-07 V_low
+ 4.412000000e-07 V_low
+ 4.412010000e-07 V_low
+ 4.413000000e-07 V_low
+ 4.413010000e-07 V_low
+ 4.414000000e-07 V_low
+ 4.414010000e-07 V_low
+ 4.415000000e-07 V_low
+ 4.415010000e-07 V_low
+ 4.416000000e-07 V_low
+ 4.416010000e-07 V_low
+ 4.417000000e-07 V_low
+ 4.417010000e-07 V_low
+ 4.418000000e-07 V_low
+ 4.418010000e-07 V_low
+ 4.419000000e-07 V_low
+ 4.419010000e-07 V_low
+ 4.420000000e-07 V_low
+ 4.420010000e-07 V_low
+ 4.421000000e-07 V_low
+ 4.421010000e-07 V_low
+ 4.422000000e-07 V_low
+ 4.422010000e-07 V_low
+ 4.423000000e-07 V_low
+ 4.423010000e-07 V_low
+ 4.424000000e-07 V_low
+ 4.424010000e-07 V_low
+ 4.425000000e-07 V_low
+ 4.425010000e-07 V_low
+ 4.426000000e-07 V_low
+ 4.426010000e-07 V_low
+ 4.427000000e-07 V_low
+ 4.427010000e-07 V_low
+ 4.428000000e-07 V_low
+ 4.428010000e-07 V_low
+ 4.429000000e-07 V_low
+ 4.429010000e-07 V_hig
+ 4.430000000e-07 V_hig
+ 4.430010000e-07 V_hig
+ 4.431000000e-07 V_hig
+ 4.431010000e-07 V_hig
+ 4.432000000e-07 V_hig
+ 4.432010000e-07 V_hig
+ 4.433000000e-07 V_hig
+ 4.433010000e-07 V_hig
+ 4.434000000e-07 V_hig
+ 4.434010000e-07 V_hig
+ 4.435000000e-07 V_hig
+ 4.435010000e-07 V_hig
+ 4.436000000e-07 V_hig
+ 4.436010000e-07 V_hig
+ 4.437000000e-07 V_hig
+ 4.437010000e-07 V_hig
+ 4.438000000e-07 V_hig
+ 4.438010000e-07 V_hig
+ 4.439000000e-07 V_hig
+ 4.439010000e-07 V_hig
+ 4.440000000e-07 V_hig
+ 4.440010000e-07 V_hig
+ 4.441000000e-07 V_hig
+ 4.441010000e-07 V_hig
+ 4.442000000e-07 V_hig
+ 4.442010000e-07 V_hig
+ 4.443000000e-07 V_hig
+ 4.443010000e-07 V_hig
+ 4.444000000e-07 V_hig
+ 4.444010000e-07 V_hig
+ 4.445000000e-07 V_hig
+ 4.445010000e-07 V_hig
+ 4.446000000e-07 V_hig
+ 4.446010000e-07 V_hig
+ 4.447000000e-07 V_hig
+ 4.447010000e-07 V_hig
+ 4.448000000e-07 V_hig
+ 4.448010000e-07 V_hig
+ 4.449000000e-07 V_hig
+ 4.449010000e-07 V_hig
+ 4.450000000e-07 V_hig
+ 4.450010000e-07 V_hig
+ 4.451000000e-07 V_hig
+ 4.451010000e-07 V_hig
+ 4.452000000e-07 V_hig
+ 4.452010000e-07 V_hig
+ 4.453000000e-07 V_hig
+ 4.453010000e-07 V_hig
+ 4.454000000e-07 V_hig
+ 4.454010000e-07 V_hig
+ 4.455000000e-07 V_hig
+ 4.455010000e-07 V_hig
+ 4.456000000e-07 V_hig
+ 4.456010000e-07 V_hig
+ 4.457000000e-07 V_hig
+ 4.457010000e-07 V_hig
+ 4.458000000e-07 V_hig
+ 4.458010000e-07 V_hig
+ 4.459000000e-07 V_hig
+ 4.459010000e-07 V_hig
+ 4.460000000e-07 V_hig
+ 4.460010000e-07 V_hig
+ 4.461000000e-07 V_hig
+ 4.461010000e-07 V_hig
+ 4.462000000e-07 V_hig
+ 4.462010000e-07 V_hig
+ 4.463000000e-07 V_hig
+ 4.463010000e-07 V_hig
+ 4.464000000e-07 V_hig
+ 4.464010000e-07 V_hig
+ 4.465000000e-07 V_hig
+ 4.465010000e-07 V_hig
+ 4.466000000e-07 V_hig
+ 4.466010000e-07 V_hig
+ 4.467000000e-07 V_hig
+ 4.467010000e-07 V_hig
+ 4.468000000e-07 V_hig
+ 4.468010000e-07 V_hig
+ 4.469000000e-07 V_hig
+ 4.469010000e-07 V_low
+ 4.470000000e-07 V_low
+ 4.470010000e-07 V_low
+ 4.471000000e-07 V_low
+ 4.471010000e-07 V_low
+ 4.472000000e-07 V_low
+ 4.472010000e-07 V_low
+ 4.473000000e-07 V_low
+ 4.473010000e-07 V_low
+ 4.474000000e-07 V_low
+ 4.474010000e-07 V_low
+ 4.475000000e-07 V_low
+ 4.475010000e-07 V_low
+ 4.476000000e-07 V_low
+ 4.476010000e-07 V_low
+ 4.477000000e-07 V_low
+ 4.477010000e-07 V_low
+ 4.478000000e-07 V_low
+ 4.478010000e-07 V_low
+ 4.479000000e-07 V_low
+ 4.479010000e-07 V_low
+ 4.480000000e-07 V_low
+ 4.480010000e-07 V_low
+ 4.481000000e-07 V_low
+ 4.481010000e-07 V_low
+ 4.482000000e-07 V_low
+ 4.482010000e-07 V_low
+ 4.483000000e-07 V_low
+ 4.483010000e-07 V_low
+ 4.484000000e-07 V_low
+ 4.484010000e-07 V_low
+ 4.485000000e-07 V_low
+ 4.485010000e-07 V_low
+ 4.486000000e-07 V_low
+ 4.486010000e-07 V_low
+ 4.487000000e-07 V_low
+ 4.487010000e-07 V_low
+ 4.488000000e-07 V_low
+ 4.488010000e-07 V_low
+ 4.489000000e-07 V_low
+ 4.489010000e-07 V_low
+ 4.490000000e-07 V_low
+ 4.490010000e-07 V_low
+ 4.491000000e-07 V_low
+ 4.491010000e-07 V_low
+ 4.492000000e-07 V_low
+ 4.492010000e-07 V_low
+ 4.493000000e-07 V_low
+ 4.493010000e-07 V_low
+ 4.494000000e-07 V_low
+ 4.494010000e-07 V_low
+ 4.495000000e-07 V_low
+ 4.495010000e-07 V_low
+ 4.496000000e-07 V_low
+ 4.496010000e-07 V_low
+ 4.497000000e-07 V_low
+ 4.497010000e-07 V_low
+ 4.498000000e-07 V_low
+ 4.498010000e-07 V_low
+ 4.499000000e-07 V_low
+ 4.499010000e-07 V_hig
+ 4.500000000e-07 V_hig
+ 4.500010000e-07 V_hig
+ 4.501000000e-07 V_hig
+ 4.501010000e-07 V_hig
+ 4.502000000e-07 V_hig
+ 4.502010000e-07 V_hig
+ 4.503000000e-07 V_hig
+ 4.503010000e-07 V_hig
+ 4.504000000e-07 V_hig
+ 4.504010000e-07 V_hig
+ 4.505000000e-07 V_hig
+ 4.505010000e-07 V_hig
+ 4.506000000e-07 V_hig
+ 4.506010000e-07 V_hig
+ 4.507000000e-07 V_hig
+ 4.507010000e-07 V_hig
+ 4.508000000e-07 V_hig
+ 4.508010000e-07 V_hig
+ 4.509000000e-07 V_hig
+ 4.509010000e-07 V_hig
+ 4.510000000e-07 V_hig
+ 4.510010000e-07 V_hig
+ 4.511000000e-07 V_hig
+ 4.511010000e-07 V_hig
+ 4.512000000e-07 V_hig
+ 4.512010000e-07 V_hig
+ 4.513000000e-07 V_hig
+ 4.513010000e-07 V_hig
+ 4.514000000e-07 V_hig
+ 4.514010000e-07 V_hig
+ 4.515000000e-07 V_hig
+ 4.515010000e-07 V_hig
+ 4.516000000e-07 V_hig
+ 4.516010000e-07 V_hig
+ 4.517000000e-07 V_hig
+ 4.517010000e-07 V_hig
+ 4.518000000e-07 V_hig
+ 4.518010000e-07 V_hig
+ 4.519000000e-07 V_hig
+ 4.519010000e-07 V_hig
+ 4.520000000e-07 V_hig
+ 4.520010000e-07 V_hig
+ 4.521000000e-07 V_hig
+ 4.521010000e-07 V_hig
+ 4.522000000e-07 V_hig
+ 4.522010000e-07 V_hig
+ 4.523000000e-07 V_hig
+ 4.523010000e-07 V_hig
+ 4.524000000e-07 V_hig
+ 4.524010000e-07 V_hig
+ 4.525000000e-07 V_hig
+ 4.525010000e-07 V_hig
+ 4.526000000e-07 V_hig
+ 4.526010000e-07 V_hig
+ 4.527000000e-07 V_hig
+ 4.527010000e-07 V_hig
+ 4.528000000e-07 V_hig
+ 4.528010000e-07 V_hig
+ 4.529000000e-07 V_hig
+ 4.529010000e-07 V_hig
+ 4.530000000e-07 V_hig
+ 4.530010000e-07 V_hig
+ 4.531000000e-07 V_hig
+ 4.531010000e-07 V_hig
+ 4.532000000e-07 V_hig
+ 4.532010000e-07 V_hig
+ 4.533000000e-07 V_hig
+ 4.533010000e-07 V_hig
+ 4.534000000e-07 V_hig
+ 4.534010000e-07 V_hig
+ 4.535000000e-07 V_hig
+ 4.535010000e-07 V_hig
+ 4.536000000e-07 V_hig
+ 4.536010000e-07 V_hig
+ 4.537000000e-07 V_hig
+ 4.537010000e-07 V_hig
+ 4.538000000e-07 V_hig
+ 4.538010000e-07 V_hig
+ 4.539000000e-07 V_hig
+ 4.539010000e-07 V_hig
+ 4.540000000e-07 V_hig
+ 4.540010000e-07 V_hig
+ 4.541000000e-07 V_hig
+ 4.541010000e-07 V_hig
+ 4.542000000e-07 V_hig
+ 4.542010000e-07 V_hig
+ 4.543000000e-07 V_hig
+ 4.543010000e-07 V_hig
+ 4.544000000e-07 V_hig
+ 4.544010000e-07 V_hig
+ 4.545000000e-07 V_hig
+ 4.545010000e-07 V_hig
+ 4.546000000e-07 V_hig
+ 4.546010000e-07 V_hig
+ 4.547000000e-07 V_hig
+ 4.547010000e-07 V_hig
+ 4.548000000e-07 V_hig
+ 4.548010000e-07 V_hig
+ 4.549000000e-07 V_hig
+ 4.549010000e-07 V_low
+ 4.550000000e-07 V_low
+ 4.550010000e-07 V_low
+ 4.551000000e-07 V_low
+ 4.551010000e-07 V_low
+ 4.552000000e-07 V_low
+ 4.552010000e-07 V_low
+ 4.553000000e-07 V_low
+ 4.553010000e-07 V_low
+ 4.554000000e-07 V_low
+ 4.554010000e-07 V_low
+ 4.555000000e-07 V_low
+ 4.555010000e-07 V_low
+ 4.556000000e-07 V_low
+ 4.556010000e-07 V_low
+ 4.557000000e-07 V_low
+ 4.557010000e-07 V_low
+ 4.558000000e-07 V_low
+ 4.558010000e-07 V_low
+ 4.559000000e-07 V_low
+ 4.559010000e-07 V_low
+ 4.560000000e-07 V_low
+ 4.560010000e-07 V_low
+ 4.561000000e-07 V_low
+ 4.561010000e-07 V_low
+ 4.562000000e-07 V_low
+ 4.562010000e-07 V_low
+ 4.563000000e-07 V_low
+ 4.563010000e-07 V_low
+ 4.564000000e-07 V_low
+ 4.564010000e-07 V_low
+ 4.565000000e-07 V_low
+ 4.565010000e-07 V_low
+ 4.566000000e-07 V_low
+ 4.566010000e-07 V_low
+ 4.567000000e-07 V_low
+ 4.567010000e-07 V_low
+ 4.568000000e-07 V_low
+ 4.568010000e-07 V_low
+ 4.569000000e-07 V_low
+ 4.569010000e-07 V_hig
+ 4.570000000e-07 V_hig
+ 4.570010000e-07 V_hig
+ 4.571000000e-07 V_hig
+ 4.571010000e-07 V_hig
+ 4.572000000e-07 V_hig
+ 4.572010000e-07 V_hig
+ 4.573000000e-07 V_hig
+ 4.573010000e-07 V_hig
+ 4.574000000e-07 V_hig
+ 4.574010000e-07 V_hig
+ 4.575000000e-07 V_hig
+ 4.575010000e-07 V_hig
+ 4.576000000e-07 V_hig
+ 4.576010000e-07 V_hig
+ 4.577000000e-07 V_hig
+ 4.577010000e-07 V_hig
+ 4.578000000e-07 V_hig
+ 4.578010000e-07 V_hig
+ 4.579000000e-07 V_hig
+ 4.579010000e-07 V_hig
+ 4.580000000e-07 V_hig
+ 4.580010000e-07 V_hig
+ 4.581000000e-07 V_hig
+ 4.581010000e-07 V_hig
+ 4.582000000e-07 V_hig
+ 4.582010000e-07 V_hig
+ 4.583000000e-07 V_hig
+ 4.583010000e-07 V_hig
+ 4.584000000e-07 V_hig
+ 4.584010000e-07 V_hig
+ 4.585000000e-07 V_hig
+ 4.585010000e-07 V_hig
+ 4.586000000e-07 V_hig
+ 4.586010000e-07 V_hig
+ 4.587000000e-07 V_hig
+ 4.587010000e-07 V_hig
+ 4.588000000e-07 V_hig
+ 4.588010000e-07 V_hig
+ 4.589000000e-07 V_hig
+ 4.589010000e-07 V_hig
+ 4.590000000e-07 V_hig
+ 4.590010000e-07 V_hig
+ 4.591000000e-07 V_hig
+ 4.591010000e-07 V_hig
+ 4.592000000e-07 V_hig
+ 4.592010000e-07 V_hig
+ 4.593000000e-07 V_hig
+ 4.593010000e-07 V_hig
+ 4.594000000e-07 V_hig
+ 4.594010000e-07 V_hig
+ 4.595000000e-07 V_hig
+ 4.595010000e-07 V_hig
+ 4.596000000e-07 V_hig
+ 4.596010000e-07 V_hig
+ 4.597000000e-07 V_hig
+ 4.597010000e-07 V_hig
+ 4.598000000e-07 V_hig
+ 4.598010000e-07 V_hig
+ 4.599000000e-07 V_hig
+ 4.599010000e-07 V_low
+ 4.600000000e-07 V_low
+ 4.600010000e-07 V_low
+ 4.601000000e-07 V_low
+ 4.601010000e-07 V_low
+ 4.602000000e-07 V_low
+ 4.602010000e-07 V_low
+ 4.603000000e-07 V_low
+ 4.603010000e-07 V_low
+ 4.604000000e-07 V_low
+ 4.604010000e-07 V_low
+ 4.605000000e-07 V_low
+ 4.605010000e-07 V_low
+ 4.606000000e-07 V_low
+ 4.606010000e-07 V_low
+ 4.607000000e-07 V_low
+ 4.607010000e-07 V_low
+ 4.608000000e-07 V_low
+ 4.608010000e-07 V_low
+ 4.609000000e-07 V_low
+ 4.609010000e-07 V_hig
+ 4.610000000e-07 V_hig
+ 4.610010000e-07 V_hig
+ 4.611000000e-07 V_hig
+ 4.611010000e-07 V_hig
+ 4.612000000e-07 V_hig
+ 4.612010000e-07 V_hig
+ 4.613000000e-07 V_hig
+ 4.613010000e-07 V_hig
+ 4.614000000e-07 V_hig
+ 4.614010000e-07 V_hig
+ 4.615000000e-07 V_hig
+ 4.615010000e-07 V_hig
+ 4.616000000e-07 V_hig
+ 4.616010000e-07 V_hig
+ 4.617000000e-07 V_hig
+ 4.617010000e-07 V_hig
+ 4.618000000e-07 V_hig
+ 4.618010000e-07 V_hig
+ 4.619000000e-07 V_hig
+ 4.619010000e-07 V_low
+ 4.620000000e-07 V_low
+ 4.620010000e-07 V_low
+ 4.621000000e-07 V_low
+ 4.621010000e-07 V_low
+ 4.622000000e-07 V_low
+ 4.622010000e-07 V_low
+ 4.623000000e-07 V_low
+ 4.623010000e-07 V_low
+ 4.624000000e-07 V_low
+ 4.624010000e-07 V_low
+ 4.625000000e-07 V_low
+ 4.625010000e-07 V_low
+ 4.626000000e-07 V_low
+ 4.626010000e-07 V_low
+ 4.627000000e-07 V_low
+ 4.627010000e-07 V_low
+ 4.628000000e-07 V_low
+ 4.628010000e-07 V_low
+ 4.629000000e-07 V_low
+ 4.629010000e-07 V_hig
+ 4.630000000e-07 V_hig
+ 4.630010000e-07 V_hig
+ 4.631000000e-07 V_hig
+ 4.631010000e-07 V_hig
+ 4.632000000e-07 V_hig
+ 4.632010000e-07 V_hig
+ 4.633000000e-07 V_hig
+ 4.633010000e-07 V_hig
+ 4.634000000e-07 V_hig
+ 4.634010000e-07 V_hig
+ 4.635000000e-07 V_hig
+ 4.635010000e-07 V_hig
+ 4.636000000e-07 V_hig
+ 4.636010000e-07 V_hig
+ 4.637000000e-07 V_hig
+ 4.637010000e-07 V_hig
+ 4.638000000e-07 V_hig
+ 4.638010000e-07 V_hig
+ 4.639000000e-07 V_hig
+ 4.639010000e-07 V_hig
+ 4.640000000e-07 V_hig
+ 4.640010000e-07 V_hig
+ 4.641000000e-07 V_hig
+ 4.641010000e-07 V_hig
+ 4.642000000e-07 V_hig
+ 4.642010000e-07 V_hig
+ 4.643000000e-07 V_hig
+ 4.643010000e-07 V_hig
+ 4.644000000e-07 V_hig
+ 4.644010000e-07 V_hig
+ 4.645000000e-07 V_hig
+ 4.645010000e-07 V_hig
+ 4.646000000e-07 V_hig
+ 4.646010000e-07 V_hig
+ 4.647000000e-07 V_hig
+ 4.647010000e-07 V_hig
+ 4.648000000e-07 V_hig
+ 4.648010000e-07 V_hig
+ 4.649000000e-07 V_hig
+ 4.649010000e-07 V_low
+ 4.650000000e-07 V_low
+ 4.650010000e-07 V_low
+ 4.651000000e-07 V_low
+ 4.651010000e-07 V_low
+ 4.652000000e-07 V_low
+ 4.652010000e-07 V_low
+ 4.653000000e-07 V_low
+ 4.653010000e-07 V_low
+ 4.654000000e-07 V_low
+ 4.654010000e-07 V_low
+ 4.655000000e-07 V_low
+ 4.655010000e-07 V_low
+ 4.656000000e-07 V_low
+ 4.656010000e-07 V_low
+ 4.657000000e-07 V_low
+ 4.657010000e-07 V_low
+ 4.658000000e-07 V_low
+ 4.658010000e-07 V_low
+ 4.659000000e-07 V_low
+ 4.659010000e-07 V_hig
+ 4.660000000e-07 V_hig
+ 4.660010000e-07 V_hig
+ 4.661000000e-07 V_hig
+ 4.661010000e-07 V_hig
+ 4.662000000e-07 V_hig
+ 4.662010000e-07 V_hig
+ 4.663000000e-07 V_hig
+ 4.663010000e-07 V_hig
+ 4.664000000e-07 V_hig
+ 4.664010000e-07 V_hig
+ 4.665000000e-07 V_hig
+ 4.665010000e-07 V_hig
+ 4.666000000e-07 V_hig
+ 4.666010000e-07 V_hig
+ 4.667000000e-07 V_hig
+ 4.667010000e-07 V_hig
+ 4.668000000e-07 V_hig
+ 4.668010000e-07 V_hig
+ 4.669000000e-07 V_hig
+ 4.669010000e-07 V_hig
+ 4.670000000e-07 V_hig
+ 4.670010000e-07 V_hig
+ 4.671000000e-07 V_hig
+ 4.671010000e-07 V_hig
+ 4.672000000e-07 V_hig
+ 4.672010000e-07 V_hig
+ 4.673000000e-07 V_hig
+ 4.673010000e-07 V_hig
+ 4.674000000e-07 V_hig
+ 4.674010000e-07 V_hig
+ 4.675000000e-07 V_hig
+ 4.675010000e-07 V_hig
+ 4.676000000e-07 V_hig
+ 4.676010000e-07 V_hig
+ 4.677000000e-07 V_hig
+ 4.677010000e-07 V_hig
+ 4.678000000e-07 V_hig
+ 4.678010000e-07 V_hig
+ 4.679000000e-07 V_hig
+ 4.679010000e-07 V_low
+ 4.680000000e-07 V_low
+ 4.680010000e-07 V_low
+ 4.681000000e-07 V_low
+ 4.681010000e-07 V_low
+ 4.682000000e-07 V_low
+ 4.682010000e-07 V_low
+ 4.683000000e-07 V_low
+ 4.683010000e-07 V_low
+ 4.684000000e-07 V_low
+ 4.684010000e-07 V_low
+ 4.685000000e-07 V_low
+ 4.685010000e-07 V_low
+ 4.686000000e-07 V_low
+ 4.686010000e-07 V_low
+ 4.687000000e-07 V_low
+ 4.687010000e-07 V_low
+ 4.688000000e-07 V_low
+ 4.688010000e-07 V_low
+ 4.689000000e-07 V_low
+ 4.689010000e-07 V_hig
+ 4.690000000e-07 V_hig
+ 4.690010000e-07 V_hig
+ 4.691000000e-07 V_hig
+ 4.691010000e-07 V_hig
+ 4.692000000e-07 V_hig
+ 4.692010000e-07 V_hig
+ 4.693000000e-07 V_hig
+ 4.693010000e-07 V_hig
+ 4.694000000e-07 V_hig
+ 4.694010000e-07 V_hig
+ 4.695000000e-07 V_hig
+ 4.695010000e-07 V_hig
+ 4.696000000e-07 V_hig
+ 4.696010000e-07 V_hig
+ 4.697000000e-07 V_hig
+ 4.697010000e-07 V_hig
+ 4.698000000e-07 V_hig
+ 4.698010000e-07 V_hig
+ 4.699000000e-07 V_hig
+ 4.699010000e-07 V_low
+ 4.700000000e-07 V_low
+ 4.700010000e-07 V_low
+ 4.701000000e-07 V_low
+ 4.701010000e-07 V_low
+ 4.702000000e-07 V_low
+ 4.702010000e-07 V_low
+ 4.703000000e-07 V_low
+ 4.703010000e-07 V_low
+ 4.704000000e-07 V_low
+ 4.704010000e-07 V_low
+ 4.705000000e-07 V_low
+ 4.705010000e-07 V_low
+ 4.706000000e-07 V_low
+ 4.706010000e-07 V_low
+ 4.707000000e-07 V_low
+ 4.707010000e-07 V_low
+ 4.708000000e-07 V_low
+ 4.708010000e-07 V_low
+ 4.709000000e-07 V_low
+ 4.709010000e-07 V_low
+ 4.710000000e-07 V_low
+ 4.710010000e-07 V_low
+ 4.711000000e-07 V_low
+ 4.711010000e-07 V_low
+ 4.712000000e-07 V_low
+ 4.712010000e-07 V_low
+ 4.713000000e-07 V_low
+ 4.713010000e-07 V_low
+ 4.714000000e-07 V_low
+ 4.714010000e-07 V_low
+ 4.715000000e-07 V_low
+ 4.715010000e-07 V_low
+ 4.716000000e-07 V_low
+ 4.716010000e-07 V_low
+ 4.717000000e-07 V_low
+ 4.717010000e-07 V_low
+ 4.718000000e-07 V_low
+ 4.718010000e-07 V_low
+ 4.719000000e-07 V_low
+ 4.719010000e-07 V_low
+ 4.720000000e-07 V_low
+ 4.720010000e-07 V_low
+ 4.721000000e-07 V_low
+ 4.721010000e-07 V_low
+ 4.722000000e-07 V_low
+ 4.722010000e-07 V_low
+ 4.723000000e-07 V_low
+ 4.723010000e-07 V_low
+ 4.724000000e-07 V_low
+ 4.724010000e-07 V_low
+ 4.725000000e-07 V_low
+ 4.725010000e-07 V_low
+ 4.726000000e-07 V_low
+ 4.726010000e-07 V_low
+ 4.727000000e-07 V_low
+ 4.727010000e-07 V_low
+ 4.728000000e-07 V_low
+ 4.728010000e-07 V_low
+ 4.729000000e-07 V_low
+ 4.729010000e-07 V_hig
+ 4.730000000e-07 V_hig
+ 4.730010000e-07 V_hig
+ 4.731000000e-07 V_hig
+ 4.731010000e-07 V_hig
+ 4.732000000e-07 V_hig
+ 4.732010000e-07 V_hig
+ 4.733000000e-07 V_hig
+ 4.733010000e-07 V_hig
+ 4.734000000e-07 V_hig
+ 4.734010000e-07 V_hig
+ 4.735000000e-07 V_hig
+ 4.735010000e-07 V_hig
+ 4.736000000e-07 V_hig
+ 4.736010000e-07 V_hig
+ 4.737000000e-07 V_hig
+ 4.737010000e-07 V_hig
+ 4.738000000e-07 V_hig
+ 4.738010000e-07 V_hig
+ 4.739000000e-07 V_hig
+ 4.739010000e-07 V_low
+ 4.740000000e-07 V_low
+ 4.740010000e-07 V_low
+ 4.741000000e-07 V_low
+ 4.741010000e-07 V_low
+ 4.742000000e-07 V_low
+ 4.742010000e-07 V_low
+ 4.743000000e-07 V_low
+ 4.743010000e-07 V_low
+ 4.744000000e-07 V_low
+ 4.744010000e-07 V_low
+ 4.745000000e-07 V_low
+ 4.745010000e-07 V_low
+ 4.746000000e-07 V_low
+ 4.746010000e-07 V_low
+ 4.747000000e-07 V_low
+ 4.747010000e-07 V_low
+ 4.748000000e-07 V_low
+ 4.748010000e-07 V_low
+ 4.749000000e-07 V_low
+ 4.749010000e-07 V_low
+ 4.750000000e-07 V_low
+ 4.750010000e-07 V_low
+ 4.751000000e-07 V_low
+ 4.751010000e-07 V_low
+ 4.752000000e-07 V_low
+ 4.752010000e-07 V_low
+ 4.753000000e-07 V_low
+ 4.753010000e-07 V_low
+ 4.754000000e-07 V_low
+ 4.754010000e-07 V_low
+ 4.755000000e-07 V_low
+ 4.755010000e-07 V_low
+ 4.756000000e-07 V_low
+ 4.756010000e-07 V_low
+ 4.757000000e-07 V_low
+ 4.757010000e-07 V_low
+ 4.758000000e-07 V_low
+ 4.758010000e-07 V_low
+ 4.759000000e-07 V_low
+ 4.759010000e-07 V_hig
+ 4.760000000e-07 V_hig
+ 4.760010000e-07 V_hig
+ 4.761000000e-07 V_hig
+ 4.761010000e-07 V_hig
+ 4.762000000e-07 V_hig
+ 4.762010000e-07 V_hig
+ 4.763000000e-07 V_hig
+ 4.763010000e-07 V_hig
+ 4.764000000e-07 V_hig
+ 4.764010000e-07 V_hig
+ 4.765000000e-07 V_hig
+ 4.765010000e-07 V_hig
+ 4.766000000e-07 V_hig
+ 4.766010000e-07 V_hig
+ 4.767000000e-07 V_hig
+ 4.767010000e-07 V_hig
+ 4.768000000e-07 V_hig
+ 4.768010000e-07 V_hig
+ 4.769000000e-07 V_hig
+ 4.769010000e-07 V_low
+ 4.770000000e-07 V_low
+ 4.770010000e-07 V_low
+ 4.771000000e-07 V_low
+ 4.771010000e-07 V_low
+ 4.772000000e-07 V_low
+ 4.772010000e-07 V_low
+ 4.773000000e-07 V_low
+ 4.773010000e-07 V_low
+ 4.774000000e-07 V_low
+ 4.774010000e-07 V_low
+ 4.775000000e-07 V_low
+ 4.775010000e-07 V_low
+ 4.776000000e-07 V_low
+ 4.776010000e-07 V_low
+ 4.777000000e-07 V_low
+ 4.777010000e-07 V_low
+ 4.778000000e-07 V_low
+ 4.778010000e-07 V_low
+ 4.779000000e-07 V_low
+ 4.779010000e-07 V_low
+ 4.780000000e-07 V_low
+ 4.780010000e-07 V_low
+ 4.781000000e-07 V_low
+ 4.781010000e-07 V_low
+ 4.782000000e-07 V_low
+ 4.782010000e-07 V_low
+ 4.783000000e-07 V_low
+ 4.783010000e-07 V_low
+ 4.784000000e-07 V_low
+ 4.784010000e-07 V_low
+ 4.785000000e-07 V_low
+ 4.785010000e-07 V_low
+ 4.786000000e-07 V_low
+ 4.786010000e-07 V_low
+ 4.787000000e-07 V_low
+ 4.787010000e-07 V_low
+ 4.788000000e-07 V_low
+ 4.788010000e-07 V_low
+ 4.789000000e-07 V_low
+ 4.789010000e-07 V_low
+ 4.790000000e-07 V_low
+ 4.790010000e-07 V_low
+ 4.791000000e-07 V_low
+ 4.791010000e-07 V_low
+ 4.792000000e-07 V_low
+ 4.792010000e-07 V_low
+ 4.793000000e-07 V_low
+ 4.793010000e-07 V_low
+ 4.794000000e-07 V_low
+ 4.794010000e-07 V_low
+ 4.795000000e-07 V_low
+ 4.795010000e-07 V_low
+ 4.796000000e-07 V_low
+ 4.796010000e-07 V_low
+ 4.797000000e-07 V_low
+ 4.797010000e-07 V_low
+ 4.798000000e-07 V_low
+ 4.798010000e-07 V_low
+ 4.799000000e-07 V_low
+ 4.799010000e-07 V_low
+ 4.800000000e-07 V_low
+ 4.800010000e-07 V_low
+ 4.801000000e-07 V_low
+ 4.801010000e-07 V_low
+ 4.802000000e-07 V_low
+ 4.802010000e-07 V_low
+ 4.803000000e-07 V_low
+ 4.803010000e-07 V_low
+ 4.804000000e-07 V_low
+ 4.804010000e-07 V_low
+ 4.805000000e-07 V_low
+ 4.805010000e-07 V_low
+ 4.806000000e-07 V_low
+ 4.806010000e-07 V_low
+ 4.807000000e-07 V_low
+ 4.807010000e-07 V_low
+ 4.808000000e-07 V_low
+ 4.808010000e-07 V_low
+ 4.809000000e-07 V_low
+ 4.809010000e-07 V_hig
+ 4.810000000e-07 V_hig
+ 4.810010000e-07 V_hig
+ 4.811000000e-07 V_hig
+ 4.811010000e-07 V_hig
+ 4.812000000e-07 V_hig
+ 4.812010000e-07 V_hig
+ 4.813000000e-07 V_hig
+ 4.813010000e-07 V_hig
+ 4.814000000e-07 V_hig
+ 4.814010000e-07 V_hig
+ 4.815000000e-07 V_hig
+ 4.815010000e-07 V_hig
+ 4.816000000e-07 V_hig
+ 4.816010000e-07 V_hig
+ 4.817000000e-07 V_hig
+ 4.817010000e-07 V_hig
+ 4.818000000e-07 V_hig
+ 4.818010000e-07 V_hig
+ 4.819000000e-07 V_hig
+ 4.819010000e-07 V_low
+ 4.820000000e-07 V_low
+ 4.820010000e-07 V_low
+ 4.821000000e-07 V_low
+ 4.821010000e-07 V_low
+ 4.822000000e-07 V_low
+ 4.822010000e-07 V_low
+ 4.823000000e-07 V_low
+ 4.823010000e-07 V_low
+ 4.824000000e-07 V_low
+ 4.824010000e-07 V_low
+ 4.825000000e-07 V_low
+ 4.825010000e-07 V_low
+ 4.826000000e-07 V_low
+ 4.826010000e-07 V_low
+ 4.827000000e-07 V_low
+ 4.827010000e-07 V_low
+ 4.828000000e-07 V_low
+ 4.828010000e-07 V_low
+ 4.829000000e-07 V_low
+ 4.829010000e-07 V_hig
+ 4.830000000e-07 V_hig
+ 4.830010000e-07 V_hig
+ 4.831000000e-07 V_hig
+ 4.831010000e-07 V_hig
+ 4.832000000e-07 V_hig
+ 4.832010000e-07 V_hig
+ 4.833000000e-07 V_hig
+ 4.833010000e-07 V_hig
+ 4.834000000e-07 V_hig
+ 4.834010000e-07 V_hig
+ 4.835000000e-07 V_hig
+ 4.835010000e-07 V_hig
+ 4.836000000e-07 V_hig
+ 4.836010000e-07 V_hig
+ 4.837000000e-07 V_hig
+ 4.837010000e-07 V_hig
+ 4.838000000e-07 V_hig
+ 4.838010000e-07 V_hig
+ 4.839000000e-07 V_hig
+ 4.839010000e-07 V_hig
+ 4.840000000e-07 V_hig
+ 4.840010000e-07 V_hig
+ 4.841000000e-07 V_hig
+ 4.841010000e-07 V_hig
+ 4.842000000e-07 V_hig
+ 4.842010000e-07 V_hig
+ 4.843000000e-07 V_hig
+ 4.843010000e-07 V_hig
+ 4.844000000e-07 V_hig
+ 4.844010000e-07 V_hig
+ 4.845000000e-07 V_hig
+ 4.845010000e-07 V_hig
+ 4.846000000e-07 V_hig
+ 4.846010000e-07 V_hig
+ 4.847000000e-07 V_hig
+ 4.847010000e-07 V_hig
+ 4.848000000e-07 V_hig
+ 4.848010000e-07 V_hig
+ 4.849000000e-07 V_hig
+ 4.849010000e-07 V_hig
+ 4.850000000e-07 V_hig
+ 4.850010000e-07 V_hig
+ 4.851000000e-07 V_hig
+ 4.851010000e-07 V_hig
+ 4.852000000e-07 V_hig
+ 4.852010000e-07 V_hig
+ 4.853000000e-07 V_hig
+ 4.853010000e-07 V_hig
+ 4.854000000e-07 V_hig
+ 4.854010000e-07 V_hig
+ 4.855000000e-07 V_hig
+ 4.855010000e-07 V_hig
+ 4.856000000e-07 V_hig
+ 4.856010000e-07 V_hig
+ 4.857000000e-07 V_hig
+ 4.857010000e-07 V_hig
+ 4.858000000e-07 V_hig
+ 4.858010000e-07 V_hig
+ 4.859000000e-07 V_hig
+ 4.859010000e-07 V_low
+ 4.860000000e-07 V_low
+ 4.860010000e-07 V_low
+ 4.861000000e-07 V_low
+ 4.861010000e-07 V_low
+ 4.862000000e-07 V_low
+ 4.862010000e-07 V_low
+ 4.863000000e-07 V_low
+ 4.863010000e-07 V_low
+ 4.864000000e-07 V_low
+ 4.864010000e-07 V_low
+ 4.865000000e-07 V_low
+ 4.865010000e-07 V_low
+ 4.866000000e-07 V_low
+ 4.866010000e-07 V_low
+ 4.867000000e-07 V_low
+ 4.867010000e-07 V_low
+ 4.868000000e-07 V_low
+ 4.868010000e-07 V_low
+ 4.869000000e-07 V_low
+ 4.869010000e-07 V_hig
+ 4.870000000e-07 V_hig
+ 4.870010000e-07 V_hig
+ 4.871000000e-07 V_hig
+ 4.871010000e-07 V_hig
+ 4.872000000e-07 V_hig
+ 4.872010000e-07 V_hig
+ 4.873000000e-07 V_hig
+ 4.873010000e-07 V_hig
+ 4.874000000e-07 V_hig
+ 4.874010000e-07 V_hig
+ 4.875000000e-07 V_hig
+ 4.875010000e-07 V_hig
+ 4.876000000e-07 V_hig
+ 4.876010000e-07 V_hig
+ 4.877000000e-07 V_hig
+ 4.877010000e-07 V_hig
+ 4.878000000e-07 V_hig
+ 4.878010000e-07 V_hig
+ 4.879000000e-07 V_hig
+ 4.879010000e-07 V_low
+ 4.880000000e-07 V_low
+ 4.880010000e-07 V_low
+ 4.881000000e-07 V_low
+ 4.881010000e-07 V_low
+ 4.882000000e-07 V_low
+ 4.882010000e-07 V_low
+ 4.883000000e-07 V_low
+ 4.883010000e-07 V_low
+ 4.884000000e-07 V_low
+ 4.884010000e-07 V_low
+ 4.885000000e-07 V_low
+ 4.885010000e-07 V_low
+ 4.886000000e-07 V_low
+ 4.886010000e-07 V_low
+ 4.887000000e-07 V_low
+ 4.887010000e-07 V_low
+ 4.888000000e-07 V_low
+ 4.888010000e-07 V_low
+ 4.889000000e-07 V_low
+ 4.889010000e-07 V_hig
+ 4.890000000e-07 V_hig
+ 4.890010000e-07 V_hig
+ 4.891000000e-07 V_hig
+ 4.891010000e-07 V_hig
+ 4.892000000e-07 V_hig
+ 4.892010000e-07 V_hig
+ 4.893000000e-07 V_hig
+ 4.893010000e-07 V_hig
+ 4.894000000e-07 V_hig
+ 4.894010000e-07 V_hig
+ 4.895000000e-07 V_hig
+ 4.895010000e-07 V_hig
+ 4.896000000e-07 V_hig
+ 4.896010000e-07 V_hig
+ 4.897000000e-07 V_hig
+ 4.897010000e-07 V_hig
+ 4.898000000e-07 V_hig
+ 4.898010000e-07 V_hig
+ 4.899000000e-07 V_hig
+ 4.899010000e-07 V_low
+ 4.900000000e-07 V_low
+ 4.900010000e-07 V_low
+ 4.901000000e-07 V_low
+ 4.901010000e-07 V_low
+ 4.902000000e-07 V_low
+ 4.902010000e-07 V_low
+ 4.903000000e-07 V_low
+ 4.903010000e-07 V_low
+ 4.904000000e-07 V_low
+ 4.904010000e-07 V_low
+ 4.905000000e-07 V_low
+ 4.905010000e-07 V_low
+ 4.906000000e-07 V_low
+ 4.906010000e-07 V_low
+ 4.907000000e-07 V_low
+ 4.907010000e-07 V_low
+ 4.908000000e-07 V_low
+ 4.908010000e-07 V_low
+ 4.909000000e-07 V_low
+ 4.909010000e-07 V_hig
+ 4.910000000e-07 V_hig
+ 4.910010000e-07 V_hig
+ 4.911000000e-07 V_hig
+ 4.911010000e-07 V_hig
+ 4.912000000e-07 V_hig
+ 4.912010000e-07 V_hig
+ 4.913000000e-07 V_hig
+ 4.913010000e-07 V_hig
+ 4.914000000e-07 V_hig
+ 4.914010000e-07 V_hig
+ 4.915000000e-07 V_hig
+ 4.915010000e-07 V_hig
+ 4.916000000e-07 V_hig
+ 4.916010000e-07 V_hig
+ 4.917000000e-07 V_hig
+ 4.917010000e-07 V_hig
+ 4.918000000e-07 V_hig
+ 4.918010000e-07 V_hig
+ 4.919000000e-07 V_hig
+ 4.919010000e-07 V_low
+ 4.920000000e-07 V_low
+ 4.920010000e-07 V_low
+ 4.921000000e-07 V_low
+ 4.921010000e-07 V_low
+ 4.922000000e-07 V_low
+ 4.922010000e-07 V_low
+ 4.923000000e-07 V_low
+ 4.923010000e-07 V_low
+ 4.924000000e-07 V_low
+ 4.924010000e-07 V_low
+ 4.925000000e-07 V_low
+ 4.925010000e-07 V_low
+ 4.926000000e-07 V_low
+ 4.926010000e-07 V_low
+ 4.927000000e-07 V_low
+ 4.927010000e-07 V_low
+ 4.928000000e-07 V_low
+ 4.928010000e-07 V_low
+ 4.929000000e-07 V_low
+ 4.929010000e-07 V_low
+ 4.930000000e-07 V_low
+ 4.930010000e-07 V_low
+ 4.931000000e-07 V_low
+ 4.931010000e-07 V_low
+ 4.932000000e-07 V_low
+ 4.932010000e-07 V_low
+ 4.933000000e-07 V_low
+ 4.933010000e-07 V_low
+ 4.934000000e-07 V_low
+ 4.934010000e-07 V_low
+ 4.935000000e-07 V_low
+ 4.935010000e-07 V_low
+ 4.936000000e-07 V_low
+ 4.936010000e-07 V_low
+ 4.937000000e-07 V_low
+ 4.937010000e-07 V_low
+ 4.938000000e-07 V_low
+ 4.938010000e-07 V_low
+ 4.939000000e-07 V_low
+ 4.939010000e-07 V_low
+ 4.940000000e-07 V_low
+ 4.940010000e-07 V_low
+ 4.941000000e-07 V_low
+ 4.941010000e-07 V_low
+ 4.942000000e-07 V_low
+ 4.942010000e-07 V_low
+ 4.943000000e-07 V_low
+ 4.943010000e-07 V_low
+ 4.944000000e-07 V_low
+ 4.944010000e-07 V_low
+ 4.945000000e-07 V_low
+ 4.945010000e-07 V_low
+ 4.946000000e-07 V_low
+ 4.946010000e-07 V_low
+ 4.947000000e-07 V_low
+ 4.947010000e-07 V_low
+ 4.948000000e-07 V_low
+ 4.948010000e-07 V_low
+ 4.949000000e-07 V_low
+ 4.949010000e-07 V_hig
+ 4.950000000e-07 V_hig
+ 4.950010000e-07 V_hig
+ 4.951000000e-07 V_hig
+ 4.951010000e-07 V_hig
+ 4.952000000e-07 V_hig
+ 4.952010000e-07 V_hig
+ 4.953000000e-07 V_hig
+ 4.953010000e-07 V_hig
+ 4.954000000e-07 V_hig
+ 4.954010000e-07 V_hig
+ 4.955000000e-07 V_hig
+ 4.955010000e-07 V_hig
+ 4.956000000e-07 V_hig
+ 4.956010000e-07 V_hig
+ 4.957000000e-07 V_hig
+ 4.957010000e-07 V_hig
+ 4.958000000e-07 V_hig
+ 4.958010000e-07 V_hig
+ 4.959000000e-07 V_hig
+ 4.959010000e-07 V_low
+ 4.960000000e-07 V_low
+ 4.960010000e-07 V_low
+ 4.961000000e-07 V_low
+ 4.961010000e-07 V_low
+ 4.962000000e-07 V_low
+ 4.962010000e-07 V_low
+ 4.963000000e-07 V_low
+ 4.963010000e-07 V_low
+ 4.964000000e-07 V_low
+ 4.964010000e-07 V_low
+ 4.965000000e-07 V_low
+ 4.965010000e-07 V_low
+ 4.966000000e-07 V_low
+ 4.966010000e-07 V_low
+ 4.967000000e-07 V_low
+ 4.967010000e-07 V_low
+ 4.968000000e-07 V_low
+ 4.968010000e-07 V_low
+ 4.969000000e-07 V_low
+ 4.969010000e-07 V_hig
+ 4.970000000e-07 V_hig
+ 4.970010000e-07 V_hig
+ 4.971000000e-07 V_hig
+ 4.971010000e-07 V_hig
+ 4.972000000e-07 V_hig
+ 4.972010000e-07 V_hig
+ 4.973000000e-07 V_hig
+ 4.973010000e-07 V_hig
+ 4.974000000e-07 V_hig
+ 4.974010000e-07 V_hig
+ 4.975000000e-07 V_hig
+ 4.975010000e-07 V_hig
+ 4.976000000e-07 V_hig
+ 4.976010000e-07 V_hig
+ 4.977000000e-07 V_hig
+ 4.977010000e-07 V_hig
+ 4.978000000e-07 V_hig
+ 4.978010000e-07 V_hig
+ 4.979000000e-07 V_hig
+ 4.979010000e-07 V_hig
+ 4.980000000e-07 V_hig
+ 4.980010000e-07 V_hig
+ 4.981000000e-07 V_hig
+ 4.981010000e-07 V_hig
+ 4.982000000e-07 V_hig
+ 4.982010000e-07 V_hig
+ 4.983000000e-07 V_hig
+ 4.983010000e-07 V_hig
+ 4.984000000e-07 V_hig
+ 4.984010000e-07 V_hig
+ 4.985000000e-07 V_hig
+ 4.985010000e-07 V_hig
+ 4.986000000e-07 V_hig
+ 4.986010000e-07 V_hig
+ 4.987000000e-07 V_hig
+ 4.987010000e-07 V_hig
+ 4.988000000e-07 V_hig
+ 4.988010000e-07 V_hig
+ 4.989000000e-07 V_hig
+ 4.989010000e-07 V_low
+ 4.990000000e-07 V_low
+ 4.990010000e-07 V_low
+ 4.991000000e-07 V_low
+ 4.991010000e-07 V_low
+ 4.992000000e-07 V_low
+ 4.992010000e-07 V_low
+ 4.993000000e-07 V_low
+ 4.993010000e-07 V_low
+ 4.994000000e-07 V_low
+ 4.994010000e-07 V_low
+ 4.995000000e-07 V_low
+ 4.995010000e-07 V_low
+ 4.996000000e-07 V_low
+ 4.996010000e-07 V_low
+ 4.997000000e-07 V_low
+ 4.997010000e-07 V_low
+ 4.998000000e-07 V_low
+ 4.998010000e-07 V_low
+ 4.999000000e-07 V_low
+ 4.999010000e-07 V_low
+ 5.000000000e-07 V_low
+ 5.000010000e-07 V_low
+ 5.001000000e-07 V_low
+ 5.001010000e-07 V_low
+ 5.002000000e-07 V_low
+ 5.002010000e-07 V_low
+ 5.003000000e-07 V_low
+ 5.003010000e-07 V_low
+ 5.004000000e-07 V_low
+ 5.004010000e-07 V_low
+ 5.005000000e-07 V_low
+ 5.005010000e-07 V_low
+ 5.006000000e-07 V_low
+ 5.006010000e-07 V_low
+ 5.007000000e-07 V_low
+ 5.007010000e-07 V_low
+ 5.008000000e-07 V_low
+ 5.008010000e-07 V_low
+ 5.009000000e-07 V_low
+ 5.009010000e-07 V_hig
+ 5.010000000e-07 V_hig
+ 5.010010000e-07 V_hig
+ 5.011000000e-07 V_hig
+ 5.011010000e-07 V_hig
+ 5.012000000e-07 V_hig
+ 5.012010000e-07 V_hig
+ 5.013000000e-07 V_hig
+ 5.013010000e-07 V_hig
+ 5.014000000e-07 V_hig
+ 5.014010000e-07 V_hig
+ 5.015000000e-07 V_hig
+ 5.015010000e-07 V_hig
+ 5.016000000e-07 V_hig
+ 5.016010000e-07 V_hig
+ 5.017000000e-07 V_hig
+ 5.017010000e-07 V_hig
+ 5.018000000e-07 V_hig
+ 5.018010000e-07 V_hig
+ 5.019000000e-07 V_hig
+ 5.019010000e-07 V_hig
+ 5.020000000e-07 V_hig
+ 5.020010000e-07 V_hig
+ 5.021000000e-07 V_hig
+ 5.021010000e-07 V_hig
+ 5.022000000e-07 V_hig
+ 5.022010000e-07 V_hig
+ 5.023000000e-07 V_hig
+ 5.023010000e-07 V_hig
+ 5.024000000e-07 V_hig
+ 5.024010000e-07 V_hig
+ 5.025000000e-07 V_hig
+ 5.025010000e-07 V_hig
+ 5.026000000e-07 V_hig
+ 5.026010000e-07 V_hig
+ 5.027000000e-07 V_hig
+ 5.027010000e-07 V_hig
+ 5.028000000e-07 V_hig
+ 5.028010000e-07 V_hig
+ 5.029000000e-07 V_hig
+ 5.029010000e-07 V_hig
+ 5.030000000e-07 V_hig
+ 5.030010000e-07 V_hig
+ 5.031000000e-07 V_hig
+ 5.031010000e-07 V_hig
+ 5.032000000e-07 V_hig
+ 5.032010000e-07 V_hig
+ 5.033000000e-07 V_hig
+ 5.033010000e-07 V_hig
+ 5.034000000e-07 V_hig
+ 5.034010000e-07 V_hig
+ 5.035000000e-07 V_hig
+ 5.035010000e-07 V_hig
+ 5.036000000e-07 V_hig
+ 5.036010000e-07 V_hig
+ 5.037000000e-07 V_hig
+ 5.037010000e-07 V_hig
+ 5.038000000e-07 V_hig
+ 5.038010000e-07 V_hig
+ 5.039000000e-07 V_hig
+ 5.039010000e-07 V_hig
+ 5.040000000e-07 V_hig
+ 5.040010000e-07 V_hig
+ 5.041000000e-07 V_hig
+ 5.041010000e-07 V_hig
+ 5.042000000e-07 V_hig
+ 5.042010000e-07 V_hig
+ 5.043000000e-07 V_hig
+ 5.043010000e-07 V_hig
+ 5.044000000e-07 V_hig
+ 5.044010000e-07 V_hig
+ 5.045000000e-07 V_hig
+ 5.045010000e-07 V_hig
+ 5.046000000e-07 V_hig
+ 5.046010000e-07 V_hig
+ 5.047000000e-07 V_hig
+ 5.047010000e-07 V_hig
+ 5.048000000e-07 V_hig
+ 5.048010000e-07 V_hig
+ 5.049000000e-07 V_hig
+ 5.049010000e-07 V_low
+ 5.050000000e-07 V_low
+ 5.050010000e-07 V_low
+ 5.051000000e-07 V_low
+ 5.051010000e-07 V_low
+ 5.052000000e-07 V_low
+ 5.052010000e-07 V_low
+ 5.053000000e-07 V_low
+ 5.053010000e-07 V_low
+ 5.054000000e-07 V_low
+ 5.054010000e-07 V_low
+ 5.055000000e-07 V_low
+ 5.055010000e-07 V_low
+ 5.056000000e-07 V_low
+ 5.056010000e-07 V_low
+ 5.057000000e-07 V_low
+ 5.057010000e-07 V_low
+ 5.058000000e-07 V_low
+ 5.058010000e-07 V_low
+ 5.059000000e-07 V_low
+ 5.059010000e-07 V_low
+ 5.060000000e-07 V_low
+ 5.060010000e-07 V_low
+ 5.061000000e-07 V_low
+ 5.061010000e-07 V_low
+ 5.062000000e-07 V_low
+ 5.062010000e-07 V_low
+ 5.063000000e-07 V_low
+ 5.063010000e-07 V_low
+ 5.064000000e-07 V_low
+ 5.064010000e-07 V_low
+ 5.065000000e-07 V_low
+ 5.065010000e-07 V_low
+ 5.066000000e-07 V_low
+ 5.066010000e-07 V_low
+ 5.067000000e-07 V_low
+ 5.067010000e-07 V_low
+ 5.068000000e-07 V_low
+ 5.068010000e-07 V_low
+ 5.069000000e-07 V_low
+ 5.069010000e-07 V_low
+ 5.070000000e-07 V_low
+ 5.070010000e-07 V_low
+ 5.071000000e-07 V_low
+ 5.071010000e-07 V_low
+ 5.072000000e-07 V_low
+ 5.072010000e-07 V_low
+ 5.073000000e-07 V_low
+ 5.073010000e-07 V_low
+ 5.074000000e-07 V_low
+ 5.074010000e-07 V_low
+ 5.075000000e-07 V_low
+ 5.075010000e-07 V_low
+ 5.076000000e-07 V_low
+ 5.076010000e-07 V_low
+ 5.077000000e-07 V_low
+ 5.077010000e-07 V_low
+ 5.078000000e-07 V_low
+ 5.078010000e-07 V_low
+ 5.079000000e-07 V_low
+ 5.079010000e-07 V_hig
+ 5.080000000e-07 V_hig
+ 5.080010000e-07 V_hig
+ 5.081000000e-07 V_hig
+ 5.081010000e-07 V_hig
+ 5.082000000e-07 V_hig
+ 5.082010000e-07 V_hig
+ 5.083000000e-07 V_hig
+ 5.083010000e-07 V_hig
+ 5.084000000e-07 V_hig
+ 5.084010000e-07 V_hig
+ 5.085000000e-07 V_hig
+ 5.085010000e-07 V_hig
+ 5.086000000e-07 V_hig
+ 5.086010000e-07 V_hig
+ 5.087000000e-07 V_hig
+ 5.087010000e-07 V_hig
+ 5.088000000e-07 V_hig
+ 5.088010000e-07 V_hig
+ 5.089000000e-07 V_hig
+ 5.089010000e-07 V_hig
+ 5.090000000e-07 V_hig
+ 5.090010000e-07 V_hig
+ 5.091000000e-07 V_hig
+ 5.091010000e-07 V_hig
+ 5.092000000e-07 V_hig
+ 5.092010000e-07 V_hig
+ 5.093000000e-07 V_hig
+ 5.093010000e-07 V_hig
+ 5.094000000e-07 V_hig
+ 5.094010000e-07 V_hig
+ 5.095000000e-07 V_hig
+ 5.095010000e-07 V_hig
+ 5.096000000e-07 V_hig
+ 5.096010000e-07 V_hig
+ 5.097000000e-07 V_hig
+ 5.097010000e-07 V_hig
+ 5.098000000e-07 V_hig
+ 5.098010000e-07 V_hig
+ 5.099000000e-07 V_hig
+ 5.099010000e-07 V_hig
+ 5.100000000e-07 V_hig
+ 5.100010000e-07 V_hig
+ 5.101000000e-07 V_hig
+ 5.101010000e-07 V_hig
+ 5.102000000e-07 V_hig
+ 5.102010000e-07 V_hig
+ 5.103000000e-07 V_hig
+ 5.103010000e-07 V_hig
+ 5.104000000e-07 V_hig
+ 5.104010000e-07 V_hig
+ 5.105000000e-07 V_hig
+ 5.105010000e-07 V_hig
+ 5.106000000e-07 V_hig
+ 5.106010000e-07 V_hig
+ 5.107000000e-07 V_hig
+ 5.107010000e-07 V_hig
+ 5.108000000e-07 V_hig
+ 5.108010000e-07 V_hig
+ 5.109000000e-07 V_hig
+ 5.109010000e-07 V_low
+ 5.110000000e-07 V_low
+ 5.110010000e-07 V_low
+ 5.111000000e-07 V_low
+ 5.111010000e-07 V_low
+ 5.112000000e-07 V_low
+ 5.112010000e-07 V_low
+ 5.113000000e-07 V_low
+ 5.113010000e-07 V_low
+ 5.114000000e-07 V_low
+ 5.114010000e-07 V_low
+ 5.115000000e-07 V_low
+ 5.115010000e-07 V_low
+ 5.116000000e-07 V_low
+ 5.116010000e-07 V_low
+ 5.117000000e-07 V_low
+ 5.117010000e-07 V_low
+ 5.118000000e-07 V_low
+ 5.118010000e-07 V_low
+ 5.119000000e-07 V_low
+ 5.119010000e-07 V_hig
+ 5.120000000e-07 V_hig
+ 5.120010000e-07 V_hig
+ 5.121000000e-07 V_hig
+ 5.121010000e-07 V_hig
+ 5.122000000e-07 V_hig
+ 5.122010000e-07 V_hig
+ 5.123000000e-07 V_hig
+ 5.123010000e-07 V_hig
+ 5.124000000e-07 V_hig
+ 5.124010000e-07 V_hig
+ 5.125000000e-07 V_hig
+ 5.125010000e-07 V_hig
+ 5.126000000e-07 V_hig
+ 5.126010000e-07 V_hig
+ 5.127000000e-07 V_hig
+ 5.127010000e-07 V_hig
+ 5.128000000e-07 V_hig
+ 5.128010000e-07 V_hig
+ 5.129000000e-07 V_hig
+ 5.129010000e-07 V_low
+ 5.130000000e-07 V_low
+ 5.130010000e-07 V_low
+ 5.131000000e-07 V_low
+ 5.131010000e-07 V_low
+ 5.132000000e-07 V_low
+ 5.132010000e-07 V_low
+ 5.133000000e-07 V_low
+ 5.133010000e-07 V_low
+ 5.134000000e-07 V_low
+ 5.134010000e-07 V_low
+ 5.135000000e-07 V_low
+ 5.135010000e-07 V_low
+ 5.136000000e-07 V_low
+ 5.136010000e-07 V_low
+ 5.137000000e-07 V_low
+ 5.137010000e-07 V_low
+ 5.138000000e-07 V_low
+ 5.138010000e-07 V_low
+ 5.139000000e-07 V_low
+ 5.139010000e-07 V_hig
+ 5.140000000e-07 V_hig
+ 5.140010000e-07 V_hig
+ 5.141000000e-07 V_hig
+ 5.141010000e-07 V_hig
+ 5.142000000e-07 V_hig
+ 5.142010000e-07 V_hig
+ 5.143000000e-07 V_hig
+ 5.143010000e-07 V_hig
+ 5.144000000e-07 V_hig
+ 5.144010000e-07 V_hig
+ 5.145000000e-07 V_hig
+ 5.145010000e-07 V_hig
+ 5.146000000e-07 V_hig
+ 5.146010000e-07 V_hig
+ 5.147000000e-07 V_hig
+ 5.147010000e-07 V_hig
+ 5.148000000e-07 V_hig
+ 5.148010000e-07 V_hig
+ 5.149000000e-07 V_hig
+ 5.149010000e-07 V_hig
+ 5.150000000e-07 V_hig
+ 5.150010000e-07 V_hig
+ 5.151000000e-07 V_hig
+ 5.151010000e-07 V_hig
+ 5.152000000e-07 V_hig
+ 5.152010000e-07 V_hig
+ 5.153000000e-07 V_hig
+ 5.153010000e-07 V_hig
+ 5.154000000e-07 V_hig
+ 5.154010000e-07 V_hig
+ 5.155000000e-07 V_hig
+ 5.155010000e-07 V_hig
+ 5.156000000e-07 V_hig
+ 5.156010000e-07 V_hig
+ 5.157000000e-07 V_hig
+ 5.157010000e-07 V_hig
+ 5.158000000e-07 V_hig
+ 5.158010000e-07 V_hig
+ 5.159000000e-07 V_hig
+ 5.159010000e-07 V_hig
+ 5.160000000e-07 V_hig
+ 5.160010000e-07 V_hig
+ 5.161000000e-07 V_hig
+ 5.161010000e-07 V_hig
+ 5.162000000e-07 V_hig
+ 5.162010000e-07 V_hig
+ 5.163000000e-07 V_hig
+ 5.163010000e-07 V_hig
+ 5.164000000e-07 V_hig
+ 5.164010000e-07 V_hig
+ 5.165000000e-07 V_hig
+ 5.165010000e-07 V_hig
+ 5.166000000e-07 V_hig
+ 5.166010000e-07 V_hig
+ 5.167000000e-07 V_hig
+ 5.167010000e-07 V_hig
+ 5.168000000e-07 V_hig
+ 5.168010000e-07 V_hig
+ 5.169000000e-07 V_hig
+ 5.169010000e-07 V_hig
+ 5.170000000e-07 V_hig
+ 5.170010000e-07 V_hig
+ 5.171000000e-07 V_hig
+ 5.171010000e-07 V_hig
+ 5.172000000e-07 V_hig
+ 5.172010000e-07 V_hig
+ 5.173000000e-07 V_hig
+ 5.173010000e-07 V_hig
+ 5.174000000e-07 V_hig
+ 5.174010000e-07 V_hig
+ 5.175000000e-07 V_hig
+ 5.175010000e-07 V_hig
+ 5.176000000e-07 V_hig
+ 5.176010000e-07 V_hig
+ 5.177000000e-07 V_hig
+ 5.177010000e-07 V_hig
+ 5.178000000e-07 V_hig
+ 5.178010000e-07 V_hig
+ 5.179000000e-07 V_hig
+ 5.179010000e-07 V_hig
+ 5.180000000e-07 V_hig
+ 5.180010000e-07 V_hig
+ 5.181000000e-07 V_hig
+ 5.181010000e-07 V_hig
+ 5.182000000e-07 V_hig
+ 5.182010000e-07 V_hig
+ 5.183000000e-07 V_hig
+ 5.183010000e-07 V_hig
+ 5.184000000e-07 V_hig
+ 5.184010000e-07 V_hig
+ 5.185000000e-07 V_hig
+ 5.185010000e-07 V_hig
+ 5.186000000e-07 V_hig
+ 5.186010000e-07 V_hig
+ 5.187000000e-07 V_hig
+ 5.187010000e-07 V_hig
+ 5.188000000e-07 V_hig
+ 5.188010000e-07 V_hig
+ 5.189000000e-07 V_hig
+ 5.189010000e-07 V_hig
+ 5.190000000e-07 V_hig
+ 5.190010000e-07 V_hig
+ 5.191000000e-07 V_hig
+ 5.191010000e-07 V_hig
+ 5.192000000e-07 V_hig
+ 5.192010000e-07 V_hig
+ 5.193000000e-07 V_hig
+ 5.193010000e-07 V_hig
+ 5.194000000e-07 V_hig
+ 5.194010000e-07 V_hig
+ 5.195000000e-07 V_hig
+ 5.195010000e-07 V_hig
+ 5.196000000e-07 V_hig
+ 5.196010000e-07 V_hig
+ 5.197000000e-07 V_hig
+ 5.197010000e-07 V_hig
+ 5.198000000e-07 V_hig
+ 5.198010000e-07 V_hig
+ 5.199000000e-07 V_hig
+ 5.199010000e-07 V_hig
+ 5.200000000e-07 V_hig
+ 5.200010000e-07 V_hig
+ 5.201000000e-07 V_hig
+ 5.201010000e-07 V_hig
+ 5.202000000e-07 V_hig
+ 5.202010000e-07 V_hig
+ 5.203000000e-07 V_hig
+ 5.203010000e-07 V_hig
+ 5.204000000e-07 V_hig
+ 5.204010000e-07 V_hig
+ 5.205000000e-07 V_hig
+ 5.205010000e-07 V_hig
+ 5.206000000e-07 V_hig
+ 5.206010000e-07 V_hig
+ 5.207000000e-07 V_hig
+ 5.207010000e-07 V_hig
+ 5.208000000e-07 V_hig
+ 5.208010000e-07 V_hig
+ 5.209000000e-07 V_hig
+ 5.209010000e-07 V_hig
+ 5.210000000e-07 V_hig
+ 5.210010000e-07 V_hig
+ 5.211000000e-07 V_hig
+ 5.211010000e-07 V_hig
+ 5.212000000e-07 V_hig
+ 5.212010000e-07 V_hig
+ 5.213000000e-07 V_hig
+ 5.213010000e-07 V_hig
+ 5.214000000e-07 V_hig
+ 5.214010000e-07 V_hig
+ 5.215000000e-07 V_hig
+ 5.215010000e-07 V_hig
+ 5.216000000e-07 V_hig
+ 5.216010000e-07 V_hig
+ 5.217000000e-07 V_hig
+ 5.217010000e-07 V_hig
+ 5.218000000e-07 V_hig
+ 5.218010000e-07 V_hig
+ 5.219000000e-07 V_hig
+ 5.219010000e-07 V_hig
+ 5.220000000e-07 V_hig
+ 5.220010000e-07 V_hig
+ 5.221000000e-07 V_hig
+ 5.221010000e-07 V_hig
+ 5.222000000e-07 V_hig
+ 5.222010000e-07 V_hig
+ 5.223000000e-07 V_hig
+ 5.223010000e-07 V_hig
+ 5.224000000e-07 V_hig
+ 5.224010000e-07 V_hig
+ 5.225000000e-07 V_hig
+ 5.225010000e-07 V_hig
+ 5.226000000e-07 V_hig
+ 5.226010000e-07 V_hig
+ 5.227000000e-07 V_hig
+ 5.227010000e-07 V_hig
+ 5.228000000e-07 V_hig
+ 5.228010000e-07 V_hig
+ 5.229000000e-07 V_hig
+ 5.229010000e-07 V_low
+ 5.230000000e-07 V_low
+ 5.230010000e-07 V_low
+ 5.231000000e-07 V_low
+ 5.231010000e-07 V_low
+ 5.232000000e-07 V_low
+ 5.232010000e-07 V_low
+ 5.233000000e-07 V_low
+ 5.233010000e-07 V_low
+ 5.234000000e-07 V_low
+ 5.234010000e-07 V_low
+ 5.235000000e-07 V_low
+ 5.235010000e-07 V_low
+ 5.236000000e-07 V_low
+ 5.236010000e-07 V_low
+ 5.237000000e-07 V_low
+ 5.237010000e-07 V_low
+ 5.238000000e-07 V_low
+ 5.238010000e-07 V_low
+ 5.239000000e-07 V_low
+ 5.239010000e-07 V_low
+ 5.240000000e-07 V_low
+ 5.240010000e-07 V_low
+ 5.241000000e-07 V_low
+ 5.241010000e-07 V_low
+ 5.242000000e-07 V_low
+ 5.242010000e-07 V_low
+ 5.243000000e-07 V_low
+ 5.243010000e-07 V_low
+ 5.244000000e-07 V_low
+ 5.244010000e-07 V_low
+ 5.245000000e-07 V_low
+ 5.245010000e-07 V_low
+ 5.246000000e-07 V_low
+ 5.246010000e-07 V_low
+ 5.247000000e-07 V_low
+ 5.247010000e-07 V_low
+ 5.248000000e-07 V_low
+ 5.248010000e-07 V_low
+ 5.249000000e-07 V_low
+ 5.249010000e-07 V_hig
+ 5.250000000e-07 V_hig
+ 5.250010000e-07 V_hig
+ 5.251000000e-07 V_hig
+ 5.251010000e-07 V_hig
+ 5.252000000e-07 V_hig
+ 5.252010000e-07 V_hig
+ 5.253000000e-07 V_hig
+ 5.253010000e-07 V_hig
+ 5.254000000e-07 V_hig
+ 5.254010000e-07 V_hig
+ 5.255000000e-07 V_hig
+ 5.255010000e-07 V_hig
+ 5.256000000e-07 V_hig
+ 5.256010000e-07 V_hig
+ 5.257000000e-07 V_hig
+ 5.257010000e-07 V_hig
+ 5.258000000e-07 V_hig
+ 5.258010000e-07 V_hig
+ 5.259000000e-07 V_hig
+ 5.259010000e-07 V_hig
+ 5.260000000e-07 V_hig
+ 5.260010000e-07 V_hig
+ 5.261000000e-07 V_hig
+ 5.261010000e-07 V_hig
+ 5.262000000e-07 V_hig
+ 5.262010000e-07 V_hig
+ 5.263000000e-07 V_hig
+ 5.263010000e-07 V_hig
+ 5.264000000e-07 V_hig
+ 5.264010000e-07 V_hig
+ 5.265000000e-07 V_hig
+ 5.265010000e-07 V_hig
+ 5.266000000e-07 V_hig
+ 5.266010000e-07 V_hig
+ 5.267000000e-07 V_hig
+ 5.267010000e-07 V_hig
+ 5.268000000e-07 V_hig
+ 5.268010000e-07 V_hig
+ 5.269000000e-07 V_hig
+ 5.269010000e-07 V_hig
+ 5.270000000e-07 V_hig
+ 5.270010000e-07 V_hig
+ 5.271000000e-07 V_hig
+ 5.271010000e-07 V_hig
+ 5.272000000e-07 V_hig
+ 5.272010000e-07 V_hig
+ 5.273000000e-07 V_hig
+ 5.273010000e-07 V_hig
+ 5.274000000e-07 V_hig
+ 5.274010000e-07 V_hig
+ 5.275000000e-07 V_hig
+ 5.275010000e-07 V_hig
+ 5.276000000e-07 V_hig
+ 5.276010000e-07 V_hig
+ 5.277000000e-07 V_hig
+ 5.277010000e-07 V_hig
+ 5.278000000e-07 V_hig
+ 5.278010000e-07 V_hig
+ 5.279000000e-07 V_hig
+ 5.279010000e-07 V_low
+ 5.280000000e-07 V_low
+ 5.280010000e-07 V_low
+ 5.281000000e-07 V_low
+ 5.281010000e-07 V_low
+ 5.282000000e-07 V_low
+ 5.282010000e-07 V_low
+ 5.283000000e-07 V_low
+ 5.283010000e-07 V_low
+ 5.284000000e-07 V_low
+ 5.284010000e-07 V_low
+ 5.285000000e-07 V_low
+ 5.285010000e-07 V_low
+ 5.286000000e-07 V_low
+ 5.286010000e-07 V_low
+ 5.287000000e-07 V_low
+ 5.287010000e-07 V_low
+ 5.288000000e-07 V_low
+ 5.288010000e-07 V_low
+ 5.289000000e-07 V_low
+ 5.289010000e-07 V_low
+ 5.290000000e-07 V_low
+ 5.290010000e-07 V_low
+ 5.291000000e-07 V_low
+ 5.291010000e-07 V_low
+ 5.292000000e-07 V_low
+ 5.292010000e-07 V_low
+ 5.293000000e-07 V_low
+ 5.293010000e-07 V_low
+ 5.294000000e-07 V_low
+ 5.294010000e-07 V_low
+ 5.295000000e-07 V_low
+ 5.295010000e-07 V_low
+ 5.296000000e-07 V_low
+ 5.296010000e-07 V_low
+ 5.297000000e-07 V_low
+ 5.297010000e-07 V_low
+ 5.298000000e-07 V_low
+ 5.298010000e-07 V_low
+ 5.299000000e-07 V_low
+ 5.299010000e-07 V_low
+ 5.300000000e-07 V_low
+ 5.300010000e-07 V_low
+ 5.301000000e-07 V_low
+ 5.301010000e-07 V_low
+ 5.302000000e-07 V_low
+ 5.302010000e-07 V_low
+ 5.303000000e-07 V_low
+ 5.303010000e-07 V_low
+ 5.304000000e-07 V_low
+ 5.304010000e-07 V_low
+ 5.305000000e-07 V_low
+ 5.305010000e-07 V_low
+ 5.306000000e-07 V_low
+ 5.306010000e-07 V_low
+ 5.307000000e-07 V_low
+ 5.307010000e-07 V_low
+ 5.308000000e-07 V_low
+ 5.308010000e-07 V_low
+ 5.309000000e-07 V_low
+ 5.309010000e-07 V_low
+ 5.310000000e-07 V_low
+ 5.310010000e-07 V_low
+ 5.311000000e-07 V_low
+ 5.311010000e-07 V_low
+ 5.312000000e-07 V_low
+ 5.312010000e-07 V_low
+ 5.313000000e-07 V_low
+ 5.313010000e-07 V_low
+ 5.314000000e-07 V_low
+ 5.314010000e-07 V_low
+ 5.315000000e-07 V_low
+ 5.315010000e-07 V_low
+ 5.316000000e-07 V_low
+ 5.316010000e-07 V_low
+ 5.317000000e-07 V_low
+ 5.317010000e-07 V_low
+ 5.318000000e-07 V_low
+ 5.318010000e-07 V_low
+ 5.319000000e-07 V_low
+ 5.319010000e-07 V_low
+ 5.320000000e-07 V_low
+ 5.320010000e-07 V_low
+ 5.321000000e-07 V_low
+ 5.321010000e-07 V_low
+ 5.322000000e-07 V_low
+ 5.322010000e-07 V_low
+ 5.323000000e-07 V_low
+ 5.323010000e-07 V_low
+ 5.324000000e-07 V_low
+ 5.324010000e-07 V_low
+ 5.325000000e-07 V_low
+ 5.325010000e-07 V_low
+ 5.326000000e-07 V_low
+ 5.326010000e-07 V_low
+ 5.327000000e-07 V_low
+ 5.327010000e-07 V_low
+ 5.328000000e-07 V_low
+ 5.328010000e-07 V_low
+ 5.329000000e-07 V_low
+ 5.329010000e-07 V_low
+ 5.330000000e-07 V_low
+ 5.330010000e-07 V_low
+ 5.331000000e-07 V_low
+ 5.331010000e-07 V_low
+ 5.332000000e-07 V_low
+ 5.332010000e-07 V_low
+ 5.333000000e-07 V_low
+ 5.333010000e-07 V_low
+ 5.334000000e-07 V_low
+ 5.334010000e-07 V_low
+ 5.335000000e-07 V_low
+ 5.335010000e-07 V_low
+ 5.336000000e-07 V_low
+ 5.336010000e-07 V_low
+ 5.337000000e-07 V_low
+ 5.337010000e-07 V_low
+ 5.338000000e-07 V_low
+ 5.338010000e-07 V_low
+ 5.339000000e-07 V_low
+ 5.339010000e-07 V_hig
+ 5.340000000e-07 V_hig
+ 5.340010000e-07 V_hig
+ 5.341000000e-07 V_hig
+ 5.341010000e-07 V_hig
+ 5.342000000e-07 V_hig
+ 5.342010000e-07 V_hig
+ 5.343000000e-07 V_hig
+ 5.343010000e-07 V_hig
+ 5.344000000e-07 V_hig
+ 5.344010000e-07 V_hig
+ 5.345000000e-07 V_hig
+ 5.345010000e-07 V_hig
+ 5.346000000e-07 V_hig
+ 5.346010000e-07 V_hig
+ 5.347000000e-07 V_hig
+ 5.347010000e-07 V_hig
+ 5.348000000e-07 V_hig
+ 5.348010000e-07 V_hig
+ 5.349000000e-07 V_hig
+ 5.349010000e-07 V_low
+ 5.350000000e-07 V_low
+ 5.350010000e-07 V_low
+ 5.351000000e-07 V_low
+ 5.351010000e-07 V_low
+ 5.352000000e-07 V_low
+ 5.352010000e-07 V_low
+ 5.353000000e-07 V_low
+ 5.353010000e-07 V_low
+ 5.354000000e-07 V_low
+ 5.354010000e-07 V_low
+ 5.355000000e-07 V_low
+ 5.355010000e-07 V_low
+ 5.356000000e-07 V_low
+ 5.356010000e-07 V_low
+ 5.357000000e-07 V_low
+ 5.357010000e-07 V_low
+ 5.358000000e-07 V_low
+ 5.358010000e-07 V_low
+ 5.359000000e-07 V_low
+ 5.359010000e-07 V_hig
+ 5.360000000e-07 V_hig
+ 5.360010000e-07 V_hig
+ 5.361000000e-07 V_hig
+ 5.361010000e-07 V_hig
+ 5.362000000e-07 V_hig
+ 5.362010000e-07 V_hig
+ 5.363000000e-07 V_hig
+ 5.363010000e-07 V_hig
+ 5.364000000e-07 V_hig
+ 5.364010000e-07 V_hig
+ 5.365000000e-07 V_hig
+ 5.365010000e-07 V_hig
+ 5.366000000e-07 V_hig
+ 5.366010000e-07 V_hig
+ 5.367000000e-07 V_hig
+ 5.367010000e-07 V_hig
+ 5.368000000e-07 V_hig
+ 5.368010000e-07 V_hig
+ 5.369000000e-07 V_hig
+ 5.369010000e-07 V_hig
+ 5.370000000e-07 V_hig
+ 5.370010000e-07 V_hig
+ 5.371000000e-07 V_hig
+ 5.371010000e-07 V_hig
+ 5.372000000e-07 V_hig
+ 5.372010000e-07 V_hig
+ 5.373000000e-07 V_hig
+ 5.373010000e-07 V_hig
+ 5.374000000e-07 V_hig
+ 5.374010000e-07 V_hig
+ 5.375000000e-07 V_hig
+ 5.375010000e-07 V_hig
+ 5.376000000e-07 V_hig
+ 5.376010000e-07 V_hig
+ 5.377000000e-07 V_hig
+ 5.377010000e-07 V_hig
+ 5.378000000e-07 V_hig
+ 5.378010000e-07 V_hig
+ 5.379000000e-07 V_hig
+ 5.379010000e-07 V_low
+ 5.380000000e-07 V_low
+ 5.380010000e-07 V_low
+ 5.381000000e-07 V_low
+ 5.381010000e-07 V_low
+ 5.382000000e-07 V_low
+ 5.382010000e-07 V_low
+ 5.383000000e-07 V_low
+ 5.383010000e-07 V_low
+ 5.384000000e-07 V_low
+ 5.384010000e-07 V_low
+ 5.385000000e-07 V_low
+ 5.385010000e-07 V_low
+ 5.386000000e-07 V_low
+ 5.386010000e-07 V_low
+ 5.387000000e-07 V_low
+ 5.387010000e-07 V_low
+ 5.388000000e-07 V_low
+ 5.388010000e-07 V_low
+ 5.389000000e-07 V_low
+ 5.389010000e-07 V_low
+ 5.390000000e-07 V_low
+ 5.390010000e-07 V_low
+ 5.391000000e-07 V_low
+ 5.391010000e-07 V_low
+ 5.392000000e-07 V_low
+ 5.392010000e-07 V_low
+ 5.393000000e-07 V_low
+ 5.393010000e-07 V_low
+ 5.394000000e-07 V_low
+ 5.394010000e-07 V_low
+ 5.395000000e-07 V_low
+ 5.395010000e-07 V_low
+ 5.396000000e-07 V_low
+ 5.396010000e-07 V_low
+ 5.397000000e-07 V_low
+ 5.397010000e-07 V_low
+ 5.398000000e-07 V_low
+ 5.398010000e-07 V_low
+ 5.399000000e-07 V_low
+ 5.399010000e-07 V_low
+ 5.400000000e-07 V_low
+ 5.400010000e-07 V_low
+ 5.401000000e-07 V_low
+ 5.401010000e-07 V_low
+ 5.402000000e-07 V_low
+ 5.402010000e-07 V_low
+ 5.403000000e-07 V_low
+ 5.403010000e-07 V_low
+ 5.404000000e-07 V_low
+ 5.404010000e-07 V_low
+ 5.405000000e-07 V_low
+ 5.405010000e-07 V_low
+ 5.406000000e-07 V_low
+ 5.406010000e-07 V_low
+ 5.407000000e-07 V_low
+ 5.407010000e-07 V_low
+ 5.408000000e-07 V_low
+ 5.408010000e-07 V_low
+ 5.409000000e-07 V_low
+ 5.409010000e-07 V_low
+ 5.410000000e-07 V_low
+ 5.410010000e-07 V_low
+ 5.411000000e-07 V_low
+ 5.411010000e-07 V_low
+ 5.412000000e-07 V_low
+ 5.412010000e-07 V_low
+ 5.413000000e-07 V_low
+ 5.413010000e-07 V_low
+ 5.414000000e-07 V_low
+ 5.414010000e-07 V_low
+ 5.415000000e-07 V_low
+ 5.415010000e-07 V_low
+ 5.416000000e-07 V_low
+ 5.416010000e-07 V_low
+ 5.417000000e-07 V_low
+ 5.417010000e-07 V_low
+ 5.418000000e-07 V_low
+ 5.418010000e-07 V_low
+ 5.419000000e-07 V_low
+ 5.419010000e-07 V_hig
+ 5.420000000e-07 V_hig
+ 5.420010000e-07 V_hig
+ 5.421000000e-07 V_hig
+ 5.421010000e-07 V_hig
+ 5.422000000e-07 V_hig
+ 5.422010000e-07 V_hig
+ 5.423000000e-07 V_hig
+ 5.423010000e-07 V_hig
+ 5.424000000e-07 V_hig
+ 5.424010000e-07 V_hig
+ 5.425000000e-07 V_hig
+ 5.425010000e-07 V_hig
+ 5.426000000e-07 V_hig
+ 5.426010000e-07 V_hig
+ 5.427000000e-07 V_hig
+ 5.427010000e-07 V_hig
+ 5.428000000e-07 V_hig
+ 5.428010000e-07 V_hig
+ 5.429000000e-07 V_hig
+ 5.429010000e-07 V_low
+ 5.430000000e-07 V_low
+ 5.430010000e-07 V_low
+ 5.431000000e-07 V_low
+ 5.431010000e-07 V_low
+ 5.432000000e-07 V_low
+ 5.432010000e-07 V_low
+ 5.433000000e-07 V_low
+ 5.433010000e-07 V_low
+ 5.434000000e-07 V_low
+ 5.434010000e-07 V_low
+ 5.435000000e-07 V_low
+ 5.435010000e-07 V_low
+ 5.436000000e-07 V_low
+ 5.436010000e-07 V_low
+ 5.437000000e-07 V_low
+ 5.437010000e-07 V_low
+ 5.438000000e-07 V_low
+ 5.438010000e-07 V_low
+ 5.439000000e-07 V_low
+ 5.439010000e-07 V_low
+ 5.440000000e-07 V_low
+ 5.440010000e-07 V_low
+ 5.441000000e-07 V_low
+ 5.441010000e-07 V_low
+ 5.442000000e-07 V_low
+ 5.442010000e-07 V_low
+ 5.443000000e-07 V_low
+ 5.443010000e-07 V_low
+ 5.444000000e-07 V_low
+ 5.444010000e-07 V_low
+ 5.445000000e-07 V_low
+ 5.445010000e-07 V_low
+ 5.446000000e-07 V_low
+ 5.446010000e-07 V_low
+ 5.447000000e-07 V_low
+ 5.447010000e-07 V_low
+ 5.448000000e-07 V_low
+ 5.448010000e-07 V_low
+ 5.449000000e-07 V_low
+ 5.449010000e-07 V_low
+ 5.450000000e-07 V_low
+ 5.450010000e-07 V_low
+ 5.451000000e-07 V_low
+ 5.451010000e-07 V_low
+ 5.452000000e-07 V_low
+ 5.452010000e-07 V_low
+ 5.453000000e-07 V_low
+ 5.453010000e-07 V_low
+ 5.454000000e-07 V_low
+ 5.454010000e-07 V_low
+ 5.455000000e-07 V_low
+ 5.455010000e-07 V_low
+ 5.456000000e-07 V_low
+ 5.456010000e-07 V_low
+ 5.457000000e-07 V_low
+ 5.457010000e-07 V_low
+ 5.458000000e-07 V_low
+ 5.458010000e-07 V_low
+ 5.459000000e-07 V_low
+ 5.459010000e-07 V_hig
+ 5.460000000e-07 V_hig
+ 5.460010000e-07 V_hig
+ 5.461000000e-07 V_hig
+ 5.461010000e-07 V_hig
+ 5.462000000e-07 V_hig
+ 5.462010000e-07 V_hig
+ 5.463000000e-07 V_hig
+ 5.463010000e-07 V_hig
+ 5.464000000e-07 V_hig
+ 5.464010000e-07 V_hig
+ 5.465000000e-07 V_hig
+ 5.465010000e-07 V_hig
+ 5.466000000e-07 V_hig
+ 5.466010000e-07 V_hig
+ 5.467000000e-07 V_hig
+ 5.467010000e-07 V_hig
+ 5.468000000e-07 V_hig
+ 5.468010000e-07 V_hig
+ 5.469000000e-07 V_hig
+ 5.469010000e-07 V_low
+ 5.470000000e-07 V_low
+ 5.470010000e-07 V_low
+ 5.471000000e-07 V_low
+ 5.471010000e-07 V_low
+ 5.472000000e-07 V_low
+ 5.472010000e-07 V_low
+ 5.473000000e-07 V_low
+ 5.473010000e-07 V_low
+ 5.474000000e-07 V_low
+ 5.474010000e-07 V_low
+ 5.475000000e-07 V_low
+ 5.475010000e-07 V_low
+ 5.476000000e-07 V_low
+ 5.476010000e-07 V_low
+ 5.477000000e-07 V_low
+ 5.477010000e-07 V_low
+ 5.478000000e-07 V_low
+ 5.478010000e-07 V_low
+ 5.479000000e-07 V_low
+ 5.479010000e-07 V_hig
+ 5.480000000e-07 V_hig
+ 5.480010000e-07 V_hig
+ 5.481000000e-07 V_hig
+ 5.481010000e-07 V_hig
+ 5.482000000e-07 V_hig
+ 5.482010000e-07 V_hig
+ 5.483000000e-07 V_hig
+ 5.483010000e-07 V_hig
+ 5.484000000e-07 V_hig
+ 5.484010000e-07 V_hig
+ 5.485000000e-07 V_hig
+ 5.485010000e-07 V_hig
+ 5.486000000e-07 V_hig
+ 5.486010000e-07 V_hig
+ 5.487000000e-07 V_hig
+ 5.487010000e-07 V_hig
+ 5.488000000e-07 V_hig
+ 5.488010000e-07 V_hig
+ 5.489000000e-07 V_hig
+ 5.489010000e-07 V_low
+ 5.490000000e-07 V_low
+ 5.490010000e-07 V_low
+ 5.491000000e-07 V_low
+ 5.491010000e-07 V_low
+ 5.492000000e-07 V_low
+ 5.492010000e-07 V_low
+ 5.493000000e-07 V_low
+ 5.493010000e-07 V_low
+ 5.494000000e-07 V_low
+ 5.494010000e-07 V_low
+ 5.495000000e-07 V_low
+ 5.495010000e-07 V_low
+ 5.496000000e-07 V_low
+ 5.496010000e-07 V_low
+ 5.497000000e-07 V_low
+ 5.497010000e-07 V_low
+ 5.498000000e-07 V_low
+ 5.498010000e-07 V_low
+ 5.499000000e-07 V_low
+ 5.499010000e-07 V_low
+ 5.500000000e-07 V_low
+ 5.500010000e-07 V_low
+ 5.501000000e-07 V_low
+ 5.501010000e-07 V_low
+ 5.502000000e-07 V_low
+ 5.502010000e-07 V_low
+ 5.503000000e-07 V_low
+ 5.503010000e-07 V_low
+ 5.504000000e-07 V_low
+ 5.504010000e-07 V_low
+ 5.505000000e-07 V_low
+ 5.505010000e-07 V_low
+ 5.506000000e-07 V_low
+ 5.506010000e-07 V_low
+ 5.507000000e-07 V_low
+ 5.507010000e-07 V_low
+ 5.508000000e-07 V_low
+ 5.508010000e-07 V_low
+ 5.509000000e-07 V_low
+ 5.509010000e-07 V_hig
+ 5.510000000e-07 V_hig
+ 5.510010000e-07 V_hig
+ 5.511000000e-07 V_hig
+ 5.511010000e-07 V_hig
+ 5.512000000e-07 V_hig
+ 5.512010000e-07 V_hig
+ 5.513000000e-07 V_hig
+ 5.513010000e-07 V_hig
+ 5.514000000e-07 V_hig
+ 5.514010000e-07 V_hig
+ 5.515000000e-07 V_hig
+ 5.515010000e-07 V_hig
+ 5.516000000e-07 V_hig
+ 5.516010000e-07 V_hig
+ 5.517000000e-07 V_hig
+ 5.517010000e-07 V_hig
+ 5.518000000e-07 V_hig
+ 5.518010000e-07 V_hig
+ 5.519000000e-07 V_hig
+ 5.519010000e-07 V_hig
+ 5.520000000e-07 V_hig
+ 5.520010000e-07 V_hig
+ 5.521000000e-07 V_hig
+ 5.521010000e-07 V_hig
+ 5.522000000e-07 V_hig
+ 5.522010000e-07 V_hig
+ 5.523000000e-07 V_hig
+ 5.523010000e-07 V_hig
+ 5.524000000e-07 V_hig
+ 5.524010000e-07 V_hig
+ 5.525000000e-07 V_hig
+ 5.525010000e-07 V_hig
+ 5.526000000e-07 V_hig
+ 5.526010000e-07 V_hig
+ 5.527000000e-07 V_hig
+ 5.527010000e-07 V_hig
+ 5.528000000e-07 V_hig
+ 5.528010000e-07 V_hig
+ 5.529000000e-07 V_hig
+ 5.529010000e-07 V_low
+ 5.530000000e-07 V_low
+ 5.530010000e-07 V_low
+ 5.531000000e-07 V_low
+ 5.531010000e-07 V_low
+ 5.532000000e-07 V_low
+ 5.532010000e-07 V_low
+ 5.533000000e-07 V_low
+ 5.533010000e-07 V_low
+ 5.534000000e-07 V_low
+ 5.534010000e-07 V_low
+ 5.535000000e-07 V_low
+ 5.535010000e-07 V_low
+ 5.536000000e-07 V_low
+ 5.536010000e-07 V_low
+ 5.537000000e-07 V_low
+ 5.537010000e-07 V_low
+ 5.538000000e-07 V_low
+ 5.538010000e-07 V_low
+ 5.539000000e-07 V_low
+ 5.539010000e-07 V_hig
+ 5.540000000e-07 V_hig
+ 5.540010000e-07 V_hig
+ 5.541000000e-07 V_hig
+ 5.541010000e-07 V_hig
+ 5.542000000e-07 V_hig
+ 5.542010000e-07 V_hig
+ 5.543000000e-07 V_hig
+ 5.543010000e-07 V_hig
+ 5.544000000e-07 V_hig
+ 5.544010000e-07 V_hig
+ 5.545000000e-07 V_hig
+ 5.545010000e-07 V_hig
+ 5.546000000e-07 V_hig
+ 5.546010000e-07 V_hig
+ 5.547000000e-07 V_hig
+ 5.547010000e-07 V_hig
+ 5.548000000e-07 V_hig
+ 5.548010000e-07 V_hig
+ 5.549000000e-07 V_hig
+ 5.549010000e-07 V_low
+ 5.550000000e-07 V_low
+ 5.550010000e-07 V_low
+ 5.551000000e-07 V_low
+ 5.551010000e-07 V_low
+ 5.552000000e-07 V_low
+ 5.552010000e-07 V_low
+ 5.553000000e-07 V_low
+ 5.553010000e-07 V_low
+ 5.554000000e-07 V_low
+ 5.554010000e-07 V_low
+ 5.555000000e-07 V_low
+ 5.555010000e-07 V_low
+ 5.556000000e-07 V_low
+ 5.556010000e-07 V_low
+ 5.557000000e-07 V_low
+ 5.557010000e-07 V_low
+ 5.558000000e-07 V_low
+ 5.558010000e-07 V_low
+ 5.559000000e-07 V_low
+ 5.559010000e-07 V_low
+ 5.560000000e-07 V_low
+ 5.560010000e-07 V_low
+ 5.561000000e-07 V_low
+ 5.561010000e-07 V_low
+ 5.562000000e-07 V_low
+ 5.562010000e-07 V_low
+ 5.563000000e-07 V_low
+ 5.563010000e-07 V_low
+ 5.564000000e-07 V_low
+ 5.564010000e-07 V_low
+ 5.565000000e-07 V_low
+ 5.565010000e-07 V_low
+ 5.566000000e-07 V_low
+ 5.566010000e-07 V_low
+ 5.567000000e-07 V_low
+ 5.567010000e-07 V_low
+ 5.568000000e-07 V_low
+ 5.568010000e-07 V_low
+ 5.569000000e-07 V_low
+ 5.569010000e-07 V_low
+ 5.570000000e-07 V_low
+ 5.570010000e-07 V_low
+ 5.571000000e-07 V_low
+ 5.571010000e-07 V_low
+ 5.572000000e-07 V_low
+ 5.572010000e-07 V_low
+ 5.573000000e-07 V_low
+ 5.573010000e-07 V_low
+ 5.574000000e-07 V_low
+ 5.574010000e-07 V_low
+ 5.575000000e-07 V_low
+ 5.575010000e-07 V_low
+ 5.576000000e-07 V_low
+ 5.576010000e-07 V_low
+ 5.577000000e-07 V_low
+ 5.577010000e-07 V_low
+ 5.578000000e-07 V_low
+ 5.578010000e-07 V_low
+ 5.579000000e-07 V_low
+ 5.579010000e-07 V_low
+ 5.580000000e-07 V_low
+ 5.580010000e-07 V_low
+ 5.581000000e-07 V_low
+ 5.581010000e-07 V_low
+ 5.582000000e-07 V_low
+ 5.582010000e-07 V_low
+ 5.583000000e-07 V_low
+ 5.583010000e-07 V_low
+ 5.584000000e-07 V_low
+ 5.584010000e-07 V_low
+ 5.585000000e-07 V_low
+ 5.585010000e-07 V_low
+ 5.586000000e-07 V_low
+ 5.586010000e-07 V_low
+ 5.587000000e-07 V_low
+ 5.587010000e-07 V_low
+ 5.588000000e-07 V_low
+ 5.588010000e-07 V_low
+ 5.589000000e-07 V_low
+ 5.589010000e-07 V_hig
+ 5.590000000e-07 V_hig
+ 5.590010000e-07 V_hig
+ 5.591000000e-07 V_hig
+ 5.591010000e-07 V_hig
+ 5.592000000e-07 V_hig
+ 5.592010000e-07 V_hig
+ 5.593000000e-07 V_hig
+ 5.593010000e-07 V_hig
+ 5.594000000e-07 V_hig
+ 5.594010000e-07 V_hig
+ 5.595000000e-07 V_hig
+ 5.595010000e-07 V_hig
+ 5.596000000e-07 V_hig
+ 5.596010000e-07 V_hig
+ 5.597000000e-07 V_hig
+ 5.597010000e-07 V_hig
+ 5.598000000e-07 V_hig
+ 5.598010000e-07 V_hig
+ 5.599000000e-07 V_hig
+ 5.599010000e-07 V_hig
+ 5.600000000e-07 V_hig
+ 5.600010000e-07 V_hig
+ 5.601000000e-07 V_hig
+ 5.601010000e-07 V_hig
+ 5.602000000e-07 V_hig
+ 5.602010000e-07 V_hig
+ 5.603000000e-07 V_hig
+ 5.603010000e-07 V_hig
+ 5.604000000e-07 V_hig
+ 5.604010000e-07 V_hig
+ 5.605000000e-07 V_hig
+ 5.605010000e-07 V_hig
+ 5.606000000e-07 V_hig
+ 5.606010000e-07 V_hig
+ 5.607000000e-07 V_hig
+ 5.607010000e-07 V_hig
+ 5.608000000e-07 V_hig
+ 5.608010000e-07 V_hig
+ 5.609000000e-07 V_hig
+ 5.609010000e-07 V_low
+ 5.610000000e-07 V_low
+ 5.610010000e-07 V_low
+ 5.611000000e-07 V_low
+ 5.611010000e-07 V_low
+ 5.612000000e-07 V_low
+ 5.612010000e-07 V_low
+ 5.613000000e-07 V_low
+ 5.613010000e-07 V_low
+ 5.614000000e-07 V_low
+ 5.614010000e-07 V_low
+ 5.615000000e-07 V_low
+ 5.615010000e-07 V_low
+ 5.616000000e-07 V_low
+ 5.616010000e-07 V_low
+ 5.617000000e-07 V_low
+ 5.617010000e-07 V_low
+ 5.618000000e-07 V_low
+ 5.618010000e-07 V_low
+ 5.619000000e-07 V_low
+ 5.619010000e-07 V_hig
+ 5.620000000e-07 V_hig
+ 5.620010000e-07 V_hig
+ 5.621000000e-07 V_hig
+ 5.621010000e-07 V_hig
+ 5.622000000e-07 V_hig
+ 5.622010000e-07 V_hig
+ 5.623000000e-07 V_hig
+ 5.623010000e-07 V_hig
+ 5.624000000e-07 V_hig
+ 5.624010000e-07 V_hig
+ 5.625000000e-07 V_hig
+ 5.625010000e-07 V_hig
+ 5.626000000e-07 V_hig
+ 5.626010000e-07 V_hig
+ 5.627000000e-07 V_hig
+ 5.627010000e-07 V_hig
+ 5.628000000e-07 V_hig
+ 5.628010000e-07 V_hig
+ 5.629000000e-07 V_hig
+ 5.629010000e-07 V_low
+ 5.630000000e-07 V_low
+ 5.630010000e-07 V_low
+ 5.631000000e-07 V_low
+ 5.631010000e-07 V_low
+ 5.632000000e-07 V_low
+ 5.632010000e-07 V_low
+ 5.633000000e-07 V_low
+ 5.633010000e-07 V_low
+ 5.634000000e-07 V_low
+ 5.634010000e-07 V_low
+ 5.635000000e-07 V_low
+ 5.635010000e-07 V_low
+ 5.636000000e-07 V_low
+ 5.636010000e-07 V_low
+ 5.637000000e-07 V_low
+ 5.637010000e-07 V_low
+ 5.638000000e-07 V_low
+ 5.638010000e-07 V_low
+ 5.639000000e-07 V_low
+ 5.639010000e-07 V_hig
+ 5.640000000e-07 V_hig
+ 5.640010000e-07 V_hig
+ 5.641000000e-07 V_hig
+ 5.641010000e-07 V_hig
+ 5.642000000e-07 V_hig
+ 5.642010000e-07 V_hig
+ 5.643000000e-07 V_hig
+ 5.643010000e-07 V_hig
+ 5.644000000e-07 V_hig
+ 5.644010000e-07 V_hig
+ 5.645000000e-07 V_hig
+ 5.645010000e-07 V_hig
+ 5.646000000e-07 V_hig
+ 5.646010000e-07 V_hig
+ 5.647000000e-07 V_hig
+ 5.647010000e-07 V_hig
+ 5.648000000e-07 V_hig
+ 5.648010000e-07 V_hig
+ 5.649000000e-07 V_hig
+ 5.649010000e-07 V_low
+ 5.650000000e-07 V_low
+ 5.650010000e-07 V_low
+ 5.651000000e-07 V_low
+ 5.651010000e-07 V_low
+ 5.652000000e-07 V_low
+ 5.652010000e-07 V_low
+ 5.653000000e-07 V_low
+ 5.653010000e-07 V_low
+ 5.654000000e-07 V_low
+ 5.654010000e-07 V_low
+ 5.655000000e-07 V_low
+ 5.655010000e-07 V_low
+ 5.656000000e-07 V_low
+ 5.656010000e-07 V_low
+ 5.657000000e-07 V_low
+ 5.657010000e-07 V_low
+ 5.658000000e-07 V_low
+ 5.658010000e-07 V_low
+ 5.659000000e-07 V_low
+ 5.659010000e-07 V_low
+ 5.660000000e-07 V_low
+ 5.660010000e-07 V_low
+ 5.661000000e-07 V_low
+ 5.661010000e-07 V_low
+ 5.662000000e-07 V_low
+ 5.662010000e-07 V_low
+ 5.663000000e-07 V_low
+ 5.663010000e-07 V_low
+ 5.664000000e-07 V_low
+ 5.664010000e-07 V_low
+ 5.665000000e-07 V_low
+ 5.665010000e-07 V_low
+ 5.666000000e-07 V_low
+ 5.666010000e-07 V_low
+ 5.667000000e-07 V_low
+ 5.667010000e-07 V_low
+ 5.668000000e-07 V_low
+ 5.668010000e-07 V_low
+ 5.669000000e-07 V_low
+ 5.669010000e-07 V_hig
+ 5.670000000e-07 V_hig
+ 5.670010000e-07 V_hig
+ 5.671000000e-07 V_hig
+ 5.671010000e-07 V_hig
+ 5.672000000e-07 V_hig
+ 5.672010000e-07 V_hig
+ 5.673000000e-07 V_hig
+ 5.673010000e-07 V_hig
+ 5.674000000e-07 V_hig
+ 5.674010000e-07 V_hig
+ 5.675000000e-07 V_hig
+ 5.675010000e-07 V_hig
+ 5.676000000e-07 V_hig
+ 5.676010000e-07 V_hig
+ 5.677000000e-07 V_hig
+ 5.677010000e-07 V_hig
+ 5.678000000e-07 V_hig
+ 5.678010000e-07 V_hig
+ 5.679000000e-07 V_hig
+ 5.679010000e-07 V_low
+ 5.680000000e-07 V_low
+ 5.680010000e-07 V_low
+ 5.681000000e-07 V_low
+ 5.681010000e-07 V_low
+ 5.682000000e-07 V_low
+ 5.682010000e-07 V_low
+ 5.683000000e-07 V_low
+ 5.683010000e-07 V_low
+ 5.684000000e-07 V_low
+ 5.684010000e-07 V_low
+ 5.685000000e-07 V_low
+ 5.685010000e-07 V_low
+ 5.686000000e-07 V_low
+ 5.686010000e-07 V_low
+ 5.687000000e-07 V_low
+ 5.687010000e-07 V_low
+ 5.688000000e-07 V_low
+ 5.688010000e-07 V_low
+ 5.689000000e-07 V_low
+ 5.689010000e-07 V_hig
+ 5.690000000e-07 V_hig
+ 5.690010000e-07 V_hig
+ 5.691000000e-07 V_hig
+ 5.691010000e-07 V_hig
+ 5.692000000e-07 V_hig
+ 5.692010000e-07 V_hig
+ 5.693000000e-07 V_hig
+ 5.693010000e-07 V_hig
+ 5.694000000e-07 V_hig
+ 5.694010000e-07 V_hig
+ 5.695000000e-07 V_hig
+ 5.695010000e-07 V_hig
+ 5.696000000e-07 V_hig
+ 5.696010000e-07 V_hig
+ 5.697000000e-07 V_hig
+ 5.697010000e-07 V_hig
+ 5.698000000e-07 V_hig
+ 5.698010000e-07 V_hig
+ 5.699000000e-07 V_hig
+ 5.699010000e-07 V_low
+ 5.700000000e-07 V_low
+ 5.700010000e-07 V_low
+ 5.701000000e-07 V_low
+ 5.701010000e-07 V_low
+ 5.702000000e-07 V_low
+ 5.702010000e-07 V_low
+ 5.703000000e-07 V_low
+ 5.703010000e-07 V_low
+ 5.704000000e-07 V_low
+ 5.704010000e-07 V_low
+ 5.705000000e-07 V_low
+ 5.705010000e-07 V_low
+ 5.706000000e-07 V_low
+ 5.706010000e-07 V_low
+ 5.707000000e-07 V_low
+ 5.707010000e-07 V_low
+ 5.708000000e-07 V_low
+ 5.708010000e-07 V_low
+ 5.709000000e-07 V_low
+ 5.709010000e-07 V_low
+ 5.710000000e-07 V_low
+ 5.710010000e-07 V_low
+ 5.711000000e-07 V_low
+ 5.711010000e-07 V_low
+ 5.712000000e-07 V_low
+ 5.712010000e-07 V_low
+ 5.713000000e-07 V_low
+ 5.713010000e-07 V_low
+ 5.714000000e-07 V_low
+ 5.714010000e-07 V_low
+ 5.715000000e-07 V_low
+ 5.715010000e-07 V_low
+ 5.716000000e-07 V_low
+ 5.716010000e-07 V_low
+ 5.717000000e-07 V_low
+ 5.717010000e-07 V_low
+ 5.718000000e-07 V_low
+ 5.718010000e-07 V_low
+ 5.719000000e-07 V_low
+ 5.719010000e-07 V_low
+ 5.720000000e-07 V_low
+ 5.720010000e-07 V_low
+ 5.721000000e-07 V_low
+ 5.721010000e-07 V_low
+ 5.722000000e-07 V_low
+ 5.722010000e-07 V_low
+ 5.723000000e-07 V_low
+ 5.723010000e-07 V_low
+ 5.724000000e-07 V_low
+ 5.724010000e-07 V_low
+ 5.725000000e-07 V_low
+ 5.725010000e-07 V_low
+ 5.726000000e-07 V_low
+ 5.726010000e-07 V_low
+ 5.727000000e-07 V_low
+ 5.727010000e-07 V_low
+ 5.728000000e-07 V_low
+ 5.728010000e-07 V_low
+ 5.729000000e-07 V_low
+ 5.729010000e-07 V_low
+ 5.730000000e-07 V_low
+ 5.730010000e-07 V_low
+ 5.731000000e-07 V_low
+ 5.731010000e-07 V_low
+ 5.732000000e-07 V_low
+ 5.732010000e-07 V_low
+ 5.733000000e-07 V_low
+ 5.733010000e-07 V_low
+ 5.734000000e-07 V_low
+ 5.734010000e-07 V_low
+ 5.735000000e-07 V_low
+ 5.735010000e-07 V_low
+ 5.736000000e-07 V_low
+ 5.736010000e-07 V_low
+ 5.737000000e-07 V_low
+ 5.737010000e-07 V_low
+ 5.738000000e-07 V_low
+ 5.738010000e-07 V_low
+ 5.739000000e-07 V_low
+ 5.739010000e-07 V_hig
+ 5.740000000e-07 V_hig
+ 5.740010000e-07 V_hig
+ 5.741000000e-07 V_hig
+ 5.741010000e-07 V_hig
+ 5.742000000e-07 V_hig
+ 5.742010000e-07 V_hig
+ 5.743000000e-07 V_hig
+ 5.743010000e-07 V_hig
+ 5.744000000e-07 V_hig
+ 5.744010000e-07 V_hig
+ 5.745000000e-07 V_hig
+ 5.745010000e-07 V_hig
+ 5.746000000e-07 V_hig
+ 5.746010000e-07 V_hig
+ 5.747000000e-07 V_hig
+ 5.747010000e-07 V_hig
+ 5.748000000e-07 V_hig
+ 5.748010000e-07 V_hig
+ 5.749000000e-07 V_hig
+ 5.749010000e-07 V_low
+ 5.750000000e-07 V_low
+ 5.750010000e-07 V_low
+ 5.751000000e-07 V_low
+ 5.751010000e-07 V_low
+ 5.752000000e-07 V_low
+ 5.752010000e-07 V_low
+ 5.753000000e-07 V_low
+ 5.753010000e-07 V_low
+ 5.754000000e-07 V_low
+ 5.754010000e-07 V_low
+ 5.755000000e-07 V_low
+ 5.755010000e-07 V_low
+ 5.756000000e-07 V_low
+ 5.756010000e-07 V_low
+ 5.757000000e-07 V_low
+ 5.757010000e-07 V_low
+ 5.758000000e-07 V_low
+ 5.758010000e-07 V_low
+ 5.759000000e-07 V_low
+ 5.759010000e-07 V_hig
+ 5.760000000e-07 V_hig
+ 5.760010000e-07 V_hig
+ 5.761000000e-07 V_hig
+ 5.761010000e-07 V_hig
+ 5.762000000e-07 V_hig
+ 5.762010000e-07 V_hig
+ 5.763000000e-07 V_hig
+ 5.763010000e-07 V_hig
+ 5.764000000e-07 V_hig
+ 5.764010000e-07 V_hig
+ 5.765000000e-07 V_hig
+ 5.765010000e-07 V_hig
+ 5.766000000e-07 V_hig
+ 5.766010000e-07 V_hig
+ 5.767000000e-07 V_hig
+ 5.767010000e-07 V_hig
+ 5.768000000e-07 V_hig
+ 5.768010000e-07 V_hig
+ 5.769000000e-07 V_hig
+ 5.769010000e-07 V_hig
+ 5.770000000e-07 V_hig
+ 5.770010000e-07 V_hig
+ 5.771000000e-07 V_hig
+ 5.771010000e-07 V_hig
+ 5.772000000e-07 V_hig
+ 5.772010000e-07 V_hig
+ 5.773000000e-07 V_hig
+ 5.773010000e-07 V_hig
+ 5.774000000e-07 V_hig
+ 5.774010000e-07 V_hig
+ 5.775000000e-07 V_hig
+ 5.775010000e-07 V_hig
+ 5.776000000e-07 V_hig
+ 5.776010000e-07 V_hig
+ 5.777000000e-07 V_hig
+ 5.777010000e-07 V_hig
+ 5.778000000e-07 V_hig
+ 5.778010000e-07 V_hig
+ 5.779000000e-07 V_hig
+ 5.779010000e-07 V_low
+ 5.780000000e-07 V_low
+ 5.780010000e-07 V_low
+ 5.781000000e-07 V_low
+ 5.781010000e-07 V_low
+ 5.782000000e-07 V_low
+ 5.782010000e-07 V_low
+ 5.783000000e-07 V_low
+ 5.783010000e-07 V_low
+ 5.784000000e-07 V_low
+ 5.784010000e-07 V_low
+ 5.785000000e-07 V_low
+ 5.785010000e-07 V_low
+ 5.786000000e-07 V_low
+ 5.786010000e-07 V_low
+ 5.787000000e-07 V_low
+ 5.787010000e-07 V_low
+ 5.788000000e-07 V_low
+ 5.788010000e-07 V_low
+ 5.789000000e-07 V_low
+ 5.789010000e-07 V_low
+ 5.790000000e-07 V_low
+ 5.790010000e-07 V_low
+ 5.791000000e-07 V_low
+ 5.791010000e-07 V_low
+ 5.792000000e-07 V_low
+ 5.792010000e-07 V_low
+ 5.793000000e-07 V_low
+ 5.793010000e-07 V_low
+ 5.794000000e-07 V_low
+ 5.794010000e-07 V_low
+ 5.795000000e-07 V_low
+ 5.795010000e-07 V_low
+ 5.796000000e-07 V_low
+ 5.796010000e-07 V_low
+ 5.797000000e-07 V_low
+ 5.797010000e-07 V_low
+ 5.798000000e-07 V_low
+ 5.798010000e-07 V_low
+ 5.799000000e-07 V_low
+ 5.799010000e-07 V_low
+ 5.800000000e-07 V_low
+ 5.800010000e-07 V_low
+ 5.801000000e-07 V_low
+ 5.801010000e-07 V_low
+ 5.802000000e-07 V_low
+ 5.802010000e-07 V_low
+ 5.803000000e-07 V_low
+ 5.803010000e-07 V_low
+ 5.804000000e-07 V_low
+ 5.804010000e-07 V_low
+ 5.805000000e-07 V_low
+ 5.805010000e-07 V_low
+ 5.806000000e-07 V_low
+ 5.806010000e-07 V_low
+ 5.807000000e-07 V_low
+ 5.807010000e-07 V_low
+ 5.808000000e-07 V_low
+ 5.808010000e-07 V_low
+ 5.809000000e-07 V_low
+ 5.809010000e-07 V_low
+ 5.810000000e-07 V_low
+ 5.810010000e-07 V_low
+ 5.811000000e-07 V_low
+ 5.811010000e-07 V_low
+ 5.812000000e-07 V_low
+ 5.812010000e-07 V_low
+ 5.813000000e-07 V_low
+ 5.813010000e-07 V_low
+ 5.814000000e-07 V_low
+ 5.814010000e-07 V_low
+ 5.815000000e-07 V_low
+ 5.815010000e-07 V_low
+ 5.816000000e-07 V_low
+ 5.816010000e-07 V_low
+ 5.817000000e-07 V_low
+ 5.817010000e-07 V_low
+ 5.818000000e-07 V_low
+ 5.818010000e-07 V_low
+ 5.819000000e-07 V_low
+ 5.819010000e-07 V_hig
+ 5.820000000e-07 V_hig
+ 5.820010000e-07 V_hig
+ 5.821000000e-07 V_hig
+ 5.821010000e-07 V_hig
+ 5.822000000e-07 V_hig
+ 5.822010000e-07 V_hig
+ 5.823000000e-07 V_hig
+ 5.823010000e-07 V_hig
+ 5.824000000e-07 V_hig
+ 5.824010000e-07 V_hig
+ 5.825000000e-07 V_hig
+ 5.825010000e-07 V_hig
+ 5.826000000e-07 V_hig
+ 5.826010000e-07 V_hig
+ 5.827000000e-07 V_hig
+ 5.827010000e-07 V_hig
+ 5.828000000e-07 V_hig
+ 5.828010000e-07 V_hig
+ 5.829000000e-07 V_hig
+ 5.829010000e-07 V_hig
+ 5.830000000e-07 V_hig
+ 5.830010000e-07 V_hig
+ 5.831000000e-07 V_hig
+ 5.831010000e-07 V_hig
+ 5.832000000e-07 V_hig
+ 5.832010000e-07 V_hig
+ 5.833000000e-07 V_hig
+ 5.833010000e-07 V_hig
+ 5.834000000e-07 V_hig
+ 5.834010000e-07 V_hig
+ 5.835000000e-07 V_hig
+ 5.835010000e-07 V_hig
+ 5.836000000e-07 V_hig
+ 5.836010000e-07 V_hig
+ 5.837000000e-07 V_hig
+ 5.837010000e-07 V_hig
+ 5.838000000e-07 V_hig
+ 5.838010000e-07 V_hig
+ 5.839000000e-07 V_hig
+ 5.839010000e-07 V_hig
+ 5.840000000e-07 V_hig
+ 5.840010000e-07 V_hig
+ 5.841000000e-07 V_hig
+ 5.841010000e-07 V_hig
+ 5.842000000e-07 V_hig
+ 5.842010000e-07 V_hig
+ 5.843000000e-07 V_hig
+ 5.843010000e-07 V_hig
+ 5.844000000e-07 V_hig
+ 5.844010000e-07 V_hig
+ 5.845000000e-07 V_hig
+ 5.845010000e-07 V_hig
+ 5.846000000e-07 V_hig
+ 5.846010000e-07 V_hig
+ 5.847000000e-07 V_hig
+ 5.847010000e-07 V_hig
+ 5.848000000e-07 V_hig
+ 5.848010000e-07 V_hig
+ 5.849000000e-07 V_hig
+ 5.849010000e-07 V_hig
+ 5.850000000e-07 V_hig
+ 5.850010000e-07 V_hig
+ 5.851000000e-07 V_hig
+ 5.851010000e-07 V_hig
+ 5.852000000e-07 V_hig
+ 5.852010000e-07 V_hig
+ 5.853000000e-07 V_hig
+ 5.853010000e-07 V_hig
+ 5.854000000e-07 V_hig
+ 5.854010000e-07 V_hig
+ 5.855000000e-07 V_hig
+ 5.855010000e-07 V_hig
+ 5.856000000e-07 V_hig
+ 5.856010000e-07 V_hig
+ 5.857000000e-07 V_hig
+ 5.857010000e-07 V_hig
+ 5.858000000e-07 V_hig
+ 5.858010000e-07 V_hig
+ 5.859000000e-07 V_hig
+ 5.859010000e-07 V_low
+ 5.860000000e-07 V_low
+ 5.860010000e-07 V_low
+ 5.861000000e-07 V_low
+ 5.861010000e-07 V_low
+ 5.862000000e-07 V_low
+ 5.862010000e-07 V_low
+ 5.863000000e-07 V_low
+ 5.863010000e-07 V_low
+ 5.864000000e-07 V_low
+ 5.864010000e-07 V_low
+ 5.865000000e-07 V_low
+ 5.865010000e-07 V_low
+ 5.866000000e-07 V_low
+ 5.866010000e-07 V_low
+ 5.867000000e-07 V_low
+ 5.867010000e-07 V_low
+ 5.868000000e-07 V_low
+ 5.868010000e-07 V_low
+ 5.869000000e-07 V_low
+ 5.869010000e-07 V_low
+ 5.870000000e-07 V_low
+ 5.870010000e-07 V_low
+ 5.871000000e-07 V_low
+ 5.871010000e-07 V_low
+ 5.872000000e-07 V_low
+ 5.872010000e-07 V_low
+ 5.873000000e-07 V_low
+ 5.873010000e-07 V_low
+ 5.874000000e-07 V_low
+ 5.874010000e-07 V_low
+ 5.875000000e-07 V_low
+ 5.875010000e-07 V_low
+ 5.876000000e-07 V_low
+ 5.876010000e-07 V_low
+ 5.877000000e-07 V_low
+ 5.877010000e-07 V_low
+ 5.878000000e-07 V_low
+ 5.878010000e-07 V_low
+ 5.879000000e-07 V_low
+ 5.879010000e-07 V_hig
+ 5.880000000e-07 V_hig
+ 5.880010000e-07 V_hig
+ 5.881000000e-07 V_hig
+ 5.881010000e-07 V_hig
+ 5.882000000e-07 V_hig
+ 5.882010000e-07 V_hig
+ 5.883000000e-07 V_hig
+ 5.883010000e-07 V_hig
+ 5.884000000e-07 V_hig
+ 5.884010000e-07 V_hig
+ 5.885000000e-07 V_hig
+ 5.885010000e-07 V_hig
+ 5.886000000e-07 V_hig
+ 5.886010000e-07 V_hig
+ 5.887000000e-07 V_hig
+ 5.887010000e-07 V_hig
+ 5.888000000e-07 V_hig
+ 5.888010000e-07 V_hig
+ 5.889000000e-07 V_hig
+ 5.889010000e-07 V_low
+ 5.890000000e-07 V_low
+ 5.890010000e-07 V_low
+ 5.891000000e-07 V_low
+ 5.891010000e-07 V_low
+ 5.892000000e-07 V_low
+ 5.892010000e-07 V_low
+ 5.893000000e-07 V_low
+ 5.893010000e-07 V_low
+ 5.894000000e-07 V_low
+ 5.894010000e-07 V_low
+ 5.895000000e-07 V_low
+ 5.895010000e-07 V_low
+ 5.896000000e-07 V_low
+ 5.896010000e-07 V_low
+ 5.897000000e-07 V_low
+ 5.897010000e-07 V_low
+ 5.898000000e-07 V_low
+ 5.898010000e-07 V_low
+ 5.899000000e-07 V_low
+ 5.899010000e-07 V_low
+ 5.900000000e-07 V_low
+ 5.900010000e-07 V_low
+ 5.901000000e-07 V_low
+ 5.901010000e-07 V_low
+ 5.902000000e-07 V_low
+ 5.902010000e-07 V_low
+ 5.903000000e-07 V_low
+ 5.903010000e-07 V_low
+ 5.904000000e-07 V_low
+ 5.904010000e-07 V_low
+ 5.905000000e-07 V_low
+ 5.905010000e-07 V_low
+ 5.906000000e-07 V_low
+ 5.906010000e-07 V_low
+ 5.907000000e-07 V_low
+ 5.907010000e-07 V_low
+ 5.908000000e-07 V_low
+ 5.908010000e-07 V_low
+ 5.909000000e-07 V_low
+ 5.909010000e-07 V_low
+ 5.910000000e-07 V_low
+ 5.910010000e-07 V_low
+ 5.911000000e-07 V_low
+ 5.911010000e-07 V_low
+ 5.912000000e-07 V_low
+ 5.912010000e-07 V_low
+ 5.913000000e-07 V_low
+ 5.913010000e-07 V_low
+ 5.914000000e-07 V_low
+ 5.914010000e-07 V_low
+ 5.915000000e-07 V_low
+ 5.915010000e-07 V_low
+ 5.916000000e-07 V_low
+ 5.916010000e-07 V_low
+ 5.917000000e-07 V_low
+ 5.917010000e-07 V_low
+ 5.918000000e-07 V_low
+ 5.918010000e-07 V_low
+ 5.919000000e-07 V_low
+ 5.919010000e-07 V_hig
+ 5.920000000e-07 V_hig
+ 5.920010000e-07 V_hig
+ 5.921000000e-07 V_hig
+ 5.921010000e-07 V_hig
+ 5.922000000e-07 V_hig
+ 5.922010000e-07 V_hig
+ 5.923000000e-07 V_hig
+ 5.923010000e-07 V_hig
+ 5.924000000e-07 V_hig
+ 5.924010000e-07 V_hig
+ 5.925000000e-07 V_hig
+ 5.925010000e-07 V_hig
+ 5.926000000e-07 V_hig
+ 5.926010000e-07 V_hig
+ 5.927000000e-07 V_hig
+ 5.927010000e-07 V_hig
+ 5.928000000e-07 V_hig
+ 5.928010000e-07 V_hig
+ 5.929000000e-07 V_hig
+ 5.929010000e-07 V_low
+ 5.930000000e-07 V_low
+ 5.930010000e-07 V_low
+ 5.931000000e-07 V_low
+ 5.931010000e-07 V_low
+ 5.932000000e-07 V_low
+ 5.932010000e-07 V_low
+ 5.933000000e-07 V_low
+ 5.933010000e-07 V_low
+ 5.934000000e-07 V_low
+ 5.934010000e-07 V_low
+ 5.935000000e-07 V_low
+ 5.935010000e-07 V_low
+ 5.936000000e-07 V_low
+ 5.936010000e-07 V_low
+ 5.937000000e-07 V_low
+ 5.937010000e-07 V_low
+ 5.938000000e-07 V_low
+ 5.938010000e-07 V_low
+ 5.939000000e-07 V_low
+ 5.939010000e-07 V_hig
+ 5.940000000e-07 V_hig
+ 5.940010000e-07 V_hig
+ 5.941000000e-07 V_hig
+ 5.941010000e-07 V_hig
+ 5.942000000e-07 V_hig
+ 5.942010000e-07 V_hig
+ 5.943000000e-07 V_hig
+ 5.943010000e-07 V_hig
+ 5.944000000e-07 V_hig
+ 5.944010000e-07 V_hig
+ 5.945000000e-07 V_hig
+ 5.945010000e-07 V_hig
+ 5.946000000e-07 V_hig
+ 5.946010000e-07 V_hig
+ 5.947000000e-07 V_hig
+ 5.947010000e-07 V_hig
+ 5.948000000e-07 V_hig
+ 5.948010000e-07 V_hig
+ 5.949000000e-07 V_hig
+ 5.949010000e-07 V_low
+ 5.950000000e-07 V_low
+ 5.950010000e-07 V_low
+ 5.951000000e-07 V_low
+ 5.951010000e-07 V_low
+ 5.952000000e-07 V_low
+ 5.952010000e-07 V_low
+ 5.953000000e-07 V_low
+ 5.953010000e-07 V_low
+ 5.954000000e-07 V_low
+ 5.954010000e-07 V_low
+ 5.955000000e-07 V_low
+ 5.955010000e-07 V_low
+ 5.956000000e-07 V_low
+ 5.956010000e-07 V_low
+ 5.957000000e-07 V_low
+ 5.957010000e-07 V_low
+ 5.958000000e-07 V_low
+ 5.958010000e-07 V_low
+ 5.959000000e-07 V_low
+ 5.959010000e-07 V_low
+ 5.960000000e-07 V_low
+ 5.960010000e-07 V_low
+ 5.961000000e-07 V_low
+ 5.961010000e-07 V_low
+ 5.962000000e-07 V_low
+ 5.962010000e-07 V_low
+ 5.963000000e-07 V_low
+ 5.963010000e-07 V_low
+ 5.964000000e-07 V_low
+ 5.964010000e-07 V_low
+ 5.965000000e-07 V_low
+ 5.965010000e-07 V_low
+ 5.966000000e-07 V_low
+ 5.966010000e-07 V_low
+ 5.967000000e-07 V_low
+ 5.967010000e-07 V_low
+ 5.968000000e-07 V_low
+ 5.968010000e-07 V_low
+ 5.969000000e-07 V_low
+ 5.969010000e-07 V_hig
+ 5.970000000e-07 V_hig
+ 5.970010000e-07 V_hig
+ 5.971000000e-07 V_hig
+ 5.971010000e-07 V_hig
+ 5.972000000e-07 V_hig
+ 5.972010000e-07 V_hig
+ 5.973000000e-07 V_hig
+ 5.973010000e-07 V_hig
+ 5.974000000e-07 V_hig
+ 5.974010000e-07 V_hig
+ 5.975000000e-07 V_hig
+ 5.975010000e-07 V_hig
+ 5.976000000e-07 V_hig
+ 5.976010000e-07 V_hig
+ 5.977000000e-07 V_hig
+ 5.977010000e-07 V_hig
+ 5.978000000e-07 V_hig
+ 5.978010000e-07 V_hig
+ 5.979000000e-07 V_hig
+ 5.979010000e-07 V_hig
+ 5.980000000e-07 V_hig
+ 5.980010000e-07 V_hig
+ 5.981000000e-07 V_hig
+ 5.981010000e-07 V_hig
+ 5.982000000e-07 V_hig
+ 5.982010000e-07 V_hig
+ 5.983000000e-07 V_hig
+ 5.983010000e-07 V_hig
+ 5.984000000e-07 V_hig
+ 5.984010000e-07 V_hig
+ 5.985000000e-07 V_hig
+ 5.985010000e-07 V_hig
+ 5.986000000e-07 V_hig
+ 5.986010000e-07 V_hig
+ 5.987000000e-07 V_hig
+ 5.987010000e-07 V_hig
+ 5.988000000e-07 V_hig
+ 5.988010000e-07 V_hig
+ 5.989000000e-07 V_hig
+ 5.989010000e-07 V_low
+ 5.990000000e-07 V_low
+ 5.990010000e-07 V_low
+ 5.991000000e-07 V_low
+ 5.991010000e-07 V_low
+ 5.992000000e-07 V_low
+ 5.992010000e-07 V_low
+ 5.993000000e-07 V_low
+ 5.993010000e-07 V_low
+ 5.994000000e-07 V_low
+ 5.994010000e-07 V_low
+ 5.995000000e-07 V_low
+ 5.995010000e-07 V_low
+ 5.996000000e-07 V_low
+ 5.996010000e-07 V_low
+ 5.997000000e-07 V_low
+ 5.997010000e-07 V_low
+ 5.998000000e-07 V_low
+ 5.998010000e-07 V_low
+ 5.999000000e-07 V_low
+ 5.999010000e-07 V_low
+ 6.000000000e-07 V_low
+ 6.000010000e-07 V_low
+ 6.001000000e-07 V_low
+ 6.001010000e-07 V_low
+ 6.002000000e-07 V_low
+ 6.002010000e-07 V_low
+ 6.003000000e-07 V_low
+ 6.003010000e-07 V_low
+ 6.004000000e-07 V_low
+ 6.004010000e-07 V_low
+ 6.005000000e-07 V_low
+ 6.005010000e-07 V_low
+ 6.006000000e-07 V_low
+ 6.006010000e-07 V_low
+ 6.007000000e-07 V_low
+ 6.007010000e-07 V_low
+ 6.008000000e-07 V_low
+ 6.008010000e-07 V_low
+ 6.009000000e-07 V_low
+ 6.009010000e-07 V_low
+ 6.010000000e-07 V_low
+ 6.010010000e-07 V_low
+ 6.011000000e-07 V_low
+ 6.011010000e-07 V_low
+ 6.012000000e-07 V_low
+ 6.012010000e-07 V_low
+ 6.013000000e-07 V_low
+ 6.013010000e-07 V_low
+ 6.014000000e-07 V_low
+ 6.014010000e-07 V_low
+ 6.015000000e-07 V_low
+ 6.015010000e-07 V_low
+ 6.016000000e-07 V_low
+ 6.016010000e-07 V_low
+ 6.017000000e-07 V_low
+ 6.017010000e-07 V_low
+ 6.018000000e-07 V_low
+ 6.018010000e-07 V_low
+ 6.019000000e-07 V_low
+ 6.019010000e-07 V_low
+ 6.020000000e-07 V_low
+ 6.020010000e-07 V_low
+ 6.021000000e-07 V_low
+ 6.021010000e-07 V_low
+ 6.022000000e-07 V_low
+ 6.022010000e-07 V_low
+ 6.023000000e-07 V_low
+ 6.023010000e-07 V_low
+ 6.024000000e-07 V_low
+ 6.024010000e-07 V_low
+ 6.025000000e-07 V_low
+ 6.025010000e-07 V_low
+ 6.026000000e-07 V_low
+ 6.026010000e-07 V_low
+ 6.027000000e-07 V_low
+ 6.027010000e-07 V_low
+ 6.028000000e-07 V_low
+ 6.028010000e-07 V_low
+ 6.029000000e-07 V_low
+ 6.029010000e-07 V_low
+ 6.030000000e-07 V_low
+ 6.030010000e-07 V_low
+ 6.031000000e-07 V_low
+ 6.031010000e-07 V_low
+ 6.032000000e-07 V_low
+ 6.032010000e-07 V_low
+ 6.033000000e-07 V_low
+ 6.033010000e-07 V_low
+ 6.034000000e-07 V_low
+ 6.034010000e-07 V_low
+ 6.035000000e-07 V_low
+ 6.035010000e-07 V_low
+ 6.036000000e-07 V_low
+ 6.036010000e-07 V_low
+ 6.037000000e-07 V_low
+ 6.037010000e-07 V_low
+ 6.038000000e-07 V_low
+ 6.038010000e-07 V_low
+ 6.039000000e-07 V_low
+ 6.039010000e-07 V_low
+ 6.040000000e-07 V_low
+ 6.040010000e-07 V_low
+ 6.041000000e-07 V_low
+ 6.041010000e-07 V_low
+ 6.042000000e-07 V_low
+ 6.042010000e-07 V_low
+ 6.043000000e-07 V_low
+ 6.043010000e-07 V_low
+ 6.044000000e-07 V_low
+ 6.044010000e-07 V_low
+ 6.045000000e-07 V_low
+ 6.045010000e-07 V_low
+ 6.046000000e-07 V_low
+ 6.046010000e-07 V_low
+ 6.047000000e-07 V_low
+ 6.047010000e-07 V_low
+ 6.048000000e-07 V_low
+ 6.048010000e-07 V_low
+ 6.049000000e-07 V_low
+ 6.049010000e-07 V_low
+ 6.050000000e-07 V_low
+ 6.050010000e-07 V_low
+ 6.051000000e-07 V_low
+ 6.051010000e-07 V_low
+ 6.052000000e-07 V_low
+ 6.052010000e-07 V_low
+ 6.053000000e-07 V_low
+ 6.053010000e-07 V_low
+ 6.054000000e-07 V_low
+ 6.054010000e-07 V_low
+ 6.055000000e-07 V_low
+ 6.055010000e-07 V_low
+ 6.056000000e-07 V_low
+ 6.056010000e-07 V_low
+ 6.057000000e-07 V_low
+ 6.057010000e-07 V_low
+ 6.058000000e-07 V_low
+ 6.058010000e-07 V_low
+ 6.059000000e-07 V_low
+ 6.059010000e-07 V_hig
+ 6.060000000e-07 V_hig
+ 6.060010000e-07 V_hig
+ 6.061000000e-07 V_hig
+ 6.061010000e-07 V_hig
+ 6.062000000e-07 V_hig
+ 6.062010000e-07 V_hig
+ 6.063000000e-07 V_hig
+ 6.063010000e-07 V_hig
+ 6.064000000e-07 V_hig
+ 6.064010000e-07 V_hig
+ 6.065000000e-07 V_hig
+ 6.065010000e-07 V_hig
+ 6.066000000e-07 V_hig
+ 6.066010000e-07 V_hig
+ 6.067000000e-07 V_hig
+ 6.067010000e-07 V_hig
+ 6.068000000e-07 V_hig
+ 6.068010000e-07 V_hig
+ 6.069000000e-07 V_hig
+ 6.069010000e-07 V_low
+ 6.070000000e-07 V_low
+ 6.070010000e-07 V_low
+ 6.071000000e-07 V_low
+ 6.071010000e-07 V_low
+ 6.072000000e-07 V_low
+ 6.072010000e-07 V_low
+ 6.073000000e-07 V_low
+ 6.073010000e-07 V_low
+ 6.074000000e-07 V_low
+ 6.074010000e-07 V_low
+ 6.075000000e-07 V_low
+ 6.075010000e-07 V_low
+ 6.076000000e-07 V_low
+ 6.076010000e-07 V_low
+ 6.077000000e-07 V_low
+ 6.077010000e-07 V_low
+ 6.078000000e-07 V_low
+ 6.078010000e-07 V_low
+ 6.079000000e-07 V_low
+ 6.079010000e-07 V_low
+ 6.080000000e-07 V_low
+ 6.080010000e-07 V_low
+ 6.081000000e-07 V_low
+ 6.081010000e-07 V_low
+ 6.082000000e-07 V_low
+ 6.082010000e-07 V_low
+ 6.083000000e-07 V_low
+ 6.083010000e-07 V_low
+ 6.084000000e-07 V_low
+ 6.084010000e-07 V_low
+ 6.085000000e-07 V_low
+ 6.085010000e-07 V_low
+ 6.086000000e-07 V_low
+ 6.086010000e-07 V_low
+ 6.087000000e-07 V_low
+ 6.087010000e-07 V_low
+ 6.088000000e-07 V_low
+ 6.088010000e-07 V_low
+ 6.089000000e-07 V_low
+ 6.089010000e-07 V_hig
+ 6.090000000e-07 V_hig
+ 6.090010000e-07 V_hig
+ 6.091000000e-07 V_hig
+ 6.091010000e-07 V_hig
+ 6.092000000e-07 V_hig
+ 6.092010000e-07 V_hig
+ 6.093000000e-07 V_hig
+ 6.093010000e-07 V_hig
+ 6.094000000e-07 V_hig
+ 6.094010000e-07 V_hig
+ 6.095000000e-07 V_hig
+ 6.095010000e-07 V_hig
+ 6.096000000e-07 V_hig
+ 6.096010000e-07 V_hig
+ 6.097000000e-07 V_hig
+ 6.097010000e-07 V_hig
+ 6.098000000e-07 V_hig
+ 6.098010000e-07 V_hig
+ 6.099000000e-07 V_hig
+ 6.099010000e-07 V_low
+ 6.100000000e-07 V_low
+ 6.100010000e-07 V_low
+ 6.101000000e-07 V_low
+ 6.101010000e-07 V_low
+ 6.102000000e-07 V_low
+ 6.102010000e-07 V_low
+ 6.103000000e-07 V_low
+ 6.103010000e-07 V_low
+ 6.104000000e-07 V_low
+ 6.104010000e-07 V_low
+ 6.105000000e-07 V_low
+ 6.105010000e-07 V_low
+ 6.106000000e-07 V_low
+ 6.106010000e-07 V_low
+ 6.107000000e-07 V_low
+ 6.107010000e-07 V_low
+ 6.108000000e-07 V_low
+ 6.108010000e-07 V_low
+ 6.109000000e-07 V_low
+ 6.109010000e-07 V_low
+ 6.110000000e-07 V_low
+ 6.110010000e-07 V_low
+ 6.111000000e-07 V_low
+ 6.111010000e-07 V_low
+ 6.112000000e-07 V_low
+ 6.112010000e-07 V_low
+ 6.113000000e-07 V_low
+ 6.113010000e-07 V_low
+ 6.114000000e-07 V_low
+ 6.114010000e-07 V_low
+ 6.115000000e-07 V_low
+ 6.115010000e-07 V_low
+ 6.116000000e-07 V_low
+ 6.116010000e-07 V_low
+ 6.117000000e-07 V_low
+ 6.117010000e-07 V_low
+ 6.118000000e-07 V_low
+ 6.118010000e-07 V_low
+ 6.119000000e-07 V_low
+ 6.119010000e-07 V_hig
+ 6.120000000e-07 V_hig
+ 6.120010000e-07 V_hig
+ 6.121000000e-07 V_hig
+ 6.121010000e-07 V_hig
+ 6.122000000e-07 V_hig
+ 6.122010000e-07 V_hig
+ 6.123000000e-07 V_hig
+ 6.123010000e-07 V_hig
+ 6.124000000e-07 V_hig
+ 6.124010000e-07 V_hig
+ 6.125000000e-07 V_hig
+ 6.125010000e-07 V_hig
+ 6.126000000e-07 V_hig
+ 6.126010000e-07 V_hig
+ 6.127000000e-07 V_hig
+ 6.127010000e-07 V_hig
+ 6.128000000e-07 V_hig
+ 6.128010000e-07 V_hig
+ 6.129000000e-07 V_hig
+ 6.129010000e-07 V_hig
+ 6.130000000e-07 V_hig
+ 6.130010000e-07 V_hig
+ 6.131000000e-07 V_hig
+ 6.131010000e-07 V_hig
+ 6.132000000e-07 V_hig
+ 6.132010000e-07 V_hig
+ 6.133000000e-07 V_hig
+ 6.133010000e-07 V_hig
+ 6.134000000e-07 V_hig
+ 6.134010000e-07 V_hig
+ 6.135000000e-07 V_hig
+ 6.135010000e-07 V_hig
+ 6.136000000e-07 V_hig
+ 6.136010000e-07 V_hig
+ 6.137000000e-07 V_hig
+ 6.137010000e-07 V_hig
+ 6.138000000e-07 V_hig
+ 6.138010000e-07 V_hig
+ 6.139000000e-07 V_hig
+ 6.139010000e-07 V_hig
+ 6.140000000e-07 V_hig
+ 6.140010000e-07 V_hig
+ 6.141000000e-07 V_hig
+ 6.141010000e-07 V_hig
+ 6.142000000e-07 V_hig
+ 6.142010000e-07 V_hig
+ 6.143000000e-07 V_hig
+ 6.143010000e-07 V_hig
+ 6.144000000e-07 V_hig
+ 6.144010000e-07 V_hig
+ 6.145000000e-07 V_hig
+ 6.145010000e-07 V_hig
+ 6.146000000e-07 V_hig
+ 6.146010000e-07 V_hig
+ 6.147000000e-07 V_hig
+ 6.147010000e-07 V_hig
+ 6.148000000e-07 V_hig
+ 6.148010000e-07 V_hig
+ 6.149000000e-07 V_hig
+ 6.149010000e-07 V_hig
+ 6.150000000e-07 V_hig
+ 6.150010000e-07 V_hig
+ 6.151000000e-07 V_hig
+ 6.151010000e-07 V_hig
+ 6.152000000e-07 V_hig
+ 6.152010000e-07 V_hig
+ 6.153000000e-07 V_hig
+ 6.153010000e-07 V_hig
+ 6.154000000e-07 V_hig
+ 6.154010000e-07 V_hig
+ 6.155000000e-07 V_hig
+ 6.155010000e-07 V_hig
+ 6.156000000e-07 V_hig
+ 6.156010000e-07 V_hig
+ 6.157000000e-07 V_hig
+ 6.157010000e-07 V_hig
+ 6.158000000e-07 V_hig
+ 6.158010000e-07 V_hig
+ 6.159000000e-07 V_hig
+ 6.159010000e-07 V_low
+ 6.160000000e-07 V_low
+ 6.160010000e-07 V_low
+ 6.161000000e-07 V_low
+ 6.161010000e-07 V_low
+ 6.162000000e-07 V_low
+ 6.162010000e-07 V_low
+ 6.163000000e-07 V_low
+ 6.163010000e-07 V_low
+ 6.164000000e-07 V_low
+ 6.164010000e-07 V_low
+ 6.165000000e-07 V_low
+ 6.165010000e-07 V_low
+ 6.166000000e-07 V_low
+ 6.166010000e-07 V_low
+ 6.167000000e-07 V_low
+ 6.167010000e-07 V_low
+ 6.168000000e-07 V_low
+ 6.168010000e-07 V_low
+ 6.169000000e-07 V_low
+ 6.169010000e-07 V_low
+ 6.170000000e-07 V_low
+ 6.170010000e-07 V_low
+ 6.171000000e-07 V_low
+ 6.171010000e-07 V_low
+ 6.172000000e-07 V_low
+ 6.172010000e-07 V_low
+ 6.173000000e-07 V_low
+ 6.173010000e-07 V_low
+ 6.174000000e-07 V_low
+ 6.174010000e-07 V_low
+ 6.175000000e-07 V_low
+ 6.175010000e-07 V_low
+ 6.176000000e-07 V_low
+ 6.176010000e-07 V_low
+ 6.177000000e-07 V_low
+ 6.177010000e-07 V_low
+ 6.178000000e-07 V_low
+ 6.178010000e-07 V_low
+ 6.179000000e-07 V_low
+ 6.179010000e-07 V_hig
+ 6.180000000e-07 V_hig
+ 6.180010000e-07 V_hig
+ 6.181000000e-07 V_hig
+ 6.181010000e-07 V_hig
+ 6.182000000e-07 V_hig
+ 6.182010000e-07 V_hig
+ 6.183000000e-07 V_hig
+ 6.183010000e-07 V_hig
+ 6.184000000e-07 V_hig
+ 6.184010000e-07 V_hig
+ 6.185000000e-07 V_hig
+ 6.185010000e-07 V_hig
+ 6.186000000e-07 V_hig
+ 6.186010000e-07 V_hig
+ 6.187000000e-07 V_hig
+ 6.187010000e-07 V_hig
+ 6.188000000e-07 V_hig
+ 6.188010000e-07 V_hig
+ 6.189000000e-07 V_hig
+ 6.189010000e-07 V_low
+ 6.190000000e-07 V_low
+ 6.190010000e-07 V_low
+ 6.191000000e-07 V_low
+ 6.191010000e-07 V_low
+ 6.192000000e-07 V_low
+ 6.192010000e-07 V_low
+ 6.193000000e-07 V_low
+ 6.193010000e-07 V_low
+ 6.194000000e-07 V_low
+ 6.194010000e-07 V_low
+ 6.195000000e-07 V_low
+ 6.195010000e-07 V_low
+ 6.196000000e-07 V_low
+ 6.196010000e-07 V_low
+ 6.197000000e-07 V_low
+ 6.197010000e-07 V_low
+ 6.198000000e-07 V_low
+ 6.198010000e-07 V_low
+ 6.199000000e-07 V_low
+ 6.199010000e-07 V_low
+ 6.200000000e-07 V_low
+ 6.200010000e-07 V_low
+ 6.201000000e-07 V_low
+ 6.201010000e-07 V_low
+ 6.202000000e-07 V_low
+ 6.202010000e-07 V_low
+ 6.203000000e-07 V_low
+ 6.203010000e-07 V_low
+ 6.204000000e-07 V_low
+ 6.204010000e-07 V_low
+ 6.205000000e-07 V_low
+ 6.205010000e-07 V_low
+ 6.206000000e-07 V_low
+ 6.206010000e-07 V_low
+ 6.207000000e-07 V_low
+ 6.207010000e-07 V_low
+ 6.208000000e-07 V_low
+ 6.208010000e-07 V_low
+ 6.209000000e-07 V_low
+ 6.209010000e-07 V_low
+ 6.210000000e-07 V_low
+ 6.210010000e-07 V_low
+ 6.211000000e-07 V_low
+ 6.211010000e-07 V_low
+ 6.212000000e-07 V_low
+ 6.212010000e-07 V_low
+ 6.213000000e-07 V_low
+ 6.213010000e-07 V_low
+ 6.214000000e-07 V_low
+ 6.214010000e-07 V_low
+ 6.215000000e-07 V_low
+ 6.215010000e-07 V_low
+ 6.216000000e-07 V_low
+ 6.216010000e-07 V_low
+ 6.217000000e-07 V_low
+ 6.217010000e-07 V_low
+ 6.218000000e-07 V_low
+ 6.218010000e-07 V_low
+ 6.219000000e-07 V_low
+ 6.219010000e-07 V_hig
+ 6.220000000e-07 V_hig
+ 6.220010000e-07 V_hig
+ 6.221000000e-07 V_hig
+ 6.221010000e-07 V_hig
+ 6.222000000e-07 V_hig
+ 6.222010000e-07 V_hig
+ 6.223000000e-07 V_hig
+ 6.223010000e-07 V_hig
+ 6.224000000e-07 V_hig
+ 6.224010000e-07 V_hig
+ 6.225000000e-07 V_hig
+ 6.225010000e-07 V_hig
+ 6.226000000e-07 V_hig
+ 6.226010000e-07 V_hig
+ 6.227000000e-07 V_hig
+ 6.227010000e-07 V_hig
+ 6.228000000e-07 V_hig
+ 6.228010000e-07 V_hig
+ 6.229000000e-07 V_hig
+ 6.229010000e-07 V_hig
+ 6.230000000e-07 V_hig
+ 6.230010000e-07 V_hig
+ 6.231000000e-07 V_hig
+ 6.231010000e-07 V_hig
+ 6.232000000e-07 V_hig
+ 6.232010000e-07 V_hig
+ 6.233000000e-07 V_hig
+ 6.233010000e-07 V_hig
+ 6.234000000e-07 V_hig
+ 6.234010000e-07 V_hig
+ 6.235000000e-07 V_hig
+ 6.235010000e-07 V_hig
+ 6.236000000e-07 V_hig
+ 6.236010000e-07 V_hig
+ 6.237000000e-07 V_hig
+ 6.237010000e-07 V_hig
+ 6.238000000e-07 V_hig
+ 6.238010000e-07 V_hig
+ 6.239000000e-07 V_hig
+ 6.239010000e-07 V_low
+ 6.240000000e-07 V_low
+ 6.240010000e-07 V_low
+ 6.241000000e-07 V_low
+ 6.241010000e-07 V_low
+ 6.242000000e-07 V_low
+ 6.242010000e-07 V_low
+ 6.243000000e-07 V_low
+ 6.243010000e-07 V_low
+ 6.244000000e-07 V_low
+ 6.244010000e-07 V_low
+ 6.245000000e-07 V_low
+ 6.245010000e-07 V_low
+ 6.246000000e-07 V_low
+ 6.246010000e-07 V_low
+ 6.247000000e-07 V_low
+ 6.247010000e-07 V_low
+ 6.248000000e-07 V_low
+ 6.248010000e-07 V_low
+ 6.249000000e-07 V_low
+ 6.249010000e-07 V_low
+ 6.250000000e-07 V_low
+ 6.250010000e-07 V_low
+ 6.251000000e-07 V_low
+ 6.251010000e-07 V_low
+ 6.252000000e-07 V_low
+ 6.252010000e-07 V_low
+ 6.253000000e-07 V_low
+ 6.253010000e-07 V_low
+ 6.254000000e-07 V_low
+ 6.254010000e-07 V_low
+ 6.255000000e-07 V_low
+ 6.255010000e-07 V_low
+ 6.256000000e-07 V_low
+ 6.256010000e-07 V_low
+ 6.257000000e-07 V_low
+ 6.257010000e-07 V_low
+ 6.258000000e-07 V_low
+ 6.258010000e-07 V_low
+ 6.259000000e-07 V_low
+ 6.259010000e-07 V_hig
+ 6.260000000e-07 V_hig
+ 6.260010000e-07 V_hig
+ 6.261000000e-07 V_hig
+ 6.261010000e-07 V_hig
+ 6.262000000e-07 V_hig
+ 6.262010000e-07 V_hig
+ 6.263000000e-07 V_hig
+ 6.263010000e-07 V_hig
+ 6.264000000e-07 V_hig
+ 6.264010000e-07 V_hig
+ 6.265000000e-07 V_hig
+ 6.265010000e-07 V_hig
+ 6.266000000e-07 V_hig
+ 6.266010000e-07 V_hig
+ 6.267000000e-07 V_hig
+ 6.267010000e-07 V_hig
+ 6.268000000e-07 V_hig
+ 6.268010000e-07 V_hig
+ 6.269000000e-07 V_hig
+ 6.269010000e-07 V_low
+ 6.270000000e-07 V_low
+ 6.270010000e-07 V_low
+ 6.271000000e-07 V_low
+ 6.271010000e-07 V_low
+ 6.272000000e-07 V_low
+ 6.272010000e-07 V_low
+ 6.273000000e-07 V_low
+ 6.273010000e-07 V_low
+ 6.274000000e-07 V_low
+ 6.274010000e-07 V_low
+ 6.275000000e-07 V_low
+ 6.275010000e-07 V_low
+ 6.276000000e-07 V_low
+ 6.276010000e-07 V_low
+ 6.277000000e-07 V_low
+ 6.277010000e-07 V_low
+ 6.278000000e-07 V_low
+ 6.278010000e-07 V_low
+ 6.279000000e-07 V_low
+ 6.279010000e-07 V_low
+ 6.280000000e-07 V_low
+ 6.280010000e-07 V_low
+ 6.281000000e-07 V_low
+ 6.281010000e-07 V_low
+ 6.282000000e-07 V_low
+ 6.282010000e-07 V_low
+ 6.283000000e-07 V_low
+ 6.283010000e-07 V_low
+ 6.284000000e-07 V_low
+ 6.284010000e-07 V_low
+ 6.285000000e-07 V_low
+ 6.285010000e-07 V_low
+ 6.286000000e-07 V_low
+ 6.286010000e-07 V_low
+ 6.287000000e-07 V_low
+ 6.287010000e-07 V_low
+ 6.288000000e-07 V_low
+ 6.288010000e-07 V_low
+ 6.289000000e-07 V_low
+ 6.289010000e-07 V_low
+ 6.290000000e-07 V_low
+ 6.290010000e-07 V_low
+ 6.291000000e-07 V_low
+ 6.291010000e-07 V_low
+ 6.292000000e-07 V_low
+ 6.292010000e-07 V_low
+ 6.293000000e-07 V_low
+ 6.293010000e-07 V_low
+ 6.294000000e-07 V_low
+ 6.294010000e-07 V_low
+ 6.295000000e-07 V_low
+ 6.295010000e-07 V_low
+ 6.296000000e-07 V_low
+ 6.296010000e-07 V_low
+ 6.297000000e-07 V_low
+ 6.297010000e-07 V_low
+ 6.298000000e-07 V_low
+ 6.298010000e-07 V_low
+ 6.299000000e-07 V_low
+ 6.299010000e-07 V_low
+ 6.300000000e-07 V_low
+ 6.300010000e-07 V_low
+ 6.301000000e-07 V_low
+ 6.301010000e-07 V_low
+ 6.302000000e-07 V_low
+ 6.302010000e-07 V_low
+ 6.303000000e-07 V_low
+ 6.303010000e-07 V_low
+ 6.304000000e-07 V_low
+ 6.304010000e-07 V_low
+ 6.305000000e-07 V_low
+ 6.305010000e-07 V_low
+ 6.306000000e-07 V_low
+ 6.306010000e-07 V_low
+ 6.307000000e-07 V_low
+ 6.307010000e-07 V_low
+ 6.308000000e-07 V_low
+ 6.308010000e-07 V_low
+ 6.309000000e-07 V_low
+ 6.309010000e-07 V_hig
+ 6.310000000e-07 V_hig
+ 6.310010000e-07 V_hig
+ 6.311000000e-07 V_hig
+ 6.311010000e-07 V_hig
+ 6.312000000e-07 V_hig
+ 6.312010000e-07 V_hig
+ 6.313000000e-07 V_hig
+ 6.313010000e-07 V_hig
+ 6.314000000e-07 V_hig
+ 6.314010000e-07 V_hig
+ 6.315000000e-07 V_hig
+ 6.315010000e-07 V_hig
+ 6.316000000e-07 V_hig
+ 6.316010000e-07 V_hig
+ 6.317000000e-07 V_hig
+ 6.317010000e-07 V_hig
+ 6.318000000e-07 V_hig
+ 6.318010000e-07 V_hig
+ 6.319000000e-07 V_hig
+ 6.319010000e-07 V_low
+ 6.320000000e-07 V_low
+ 6.320010000e-07 V_low
+ 6.321000000e-07 V_low
+ 6.321010000e-07 V_low
+ 6.322000000e-07 V_low
+ 6.322010000e-07 V_low
+ 6.323000000e-07 V_low
+ 6.323010000e-07 V_low
+ 6.324000000e-07 V_low
+ 6.324010000e-07 V_low
+ 6.325000000e-07 V_low
+ 6.325010000e-07 V_low
+ 6.326000000e-07 V_low
+ 6.326010000e-07 V_low
+ 6.327000000e-07 V_low
+ 6.327010000e-07 V_low
+ 6.328000000e-07 V_low
+ 6.328010000e-07 V_low
+ 6.329000000e-07 V_low
+ 6.329010000e-07 V_hig
+ 6.330000000e-07 V_hig
+ 6.330010000e-07 V_hig
+ 6.331000000e-07 V_hig
+ 6.331010000e-07 V_hig
+ 6.332000000e-07 V_hig
+ 6.332010000e-07 V_hig
+ 6.333000000e-07 V_hig
+ 6.333010000e-07 V_hig
+ 6.334000000e-07 V_hig
+ 6.334010000e-07 V_hig
+ 6.335000000e-07 V_hig
+ 6.335010000e-07 V_hig
+ 6.336000000e-07 V_hig
+ 6.336010000e-07 V_hig
+ 6.337000000e-07 V_hig
+ 6.337010000e-07 V_hig
+ 6.338000000e-07 V_hig
+ 6.338010000e-07 V_hig
+ 6.339000000e-07 V_hig
+ 6.339010000e-07 V_low
+ 6.340000000e-07 V_low
+ 6.340010000e-07 V_low
+ 6.341000000e-07 V_low
+ 6.341010000e-07 V_low
+ 6.342000000e-07 V_low
+ 6.342010000e-07 V_low
+ 6.343000000e-07 V_low
+ 6.343010000e-07 V_low
+ 6.344000000e-07 V_low
+ 6.344010000e-07 V_low
+ 6.345000000e-07 V_low
+ 6.345010000e-07 V_low
+ 6.346000000e-07 V_low
+ 6.346010000e-07 V_low
+ 6.347000000e-07 V_low
+ 6.347010000e-07 V_low
+ 6.348000000e-07 V_low
+ 6.348010000e-07 V_low
+ 6.349000000e-07 V_low
+ 6.349010000e-07 V_hig
+ 6.350000000e-07 V_hig
+ 6.350010000e-07 V_hig
+ 6.351000000e-07 V_hig
+ 6.351010000e-07 V_hig
+ 6.352000000e-07 V_hig
+ 6.352010000e-07 V_hig
+ 6.353000000e-07 V_hig
+ 6.353010000e-07 V_hig
+ 6.354000000e-07 V_hig
+ 6.354010000e-07 V_hig
+ 6.355000000e-07 V_hig
+ 6.355010000e-07 V_hig
+ 6.356000000e-07 V_hig
+ 6.356010000e-07 V_hig
+ 6.357000000e-07 V_hig
+ 6.357010000e-07 V_hig
+ 6.358000000e-07 V_hig
+ 6.358010000e-07 V_hig
+ 6.359000000e-07 V_hig
+ 6.359010000e-07 V_hig
+ 6.360000000e-07 V_hig
+ 6.360010000e-07 V_hig
+ 6.361000000e-07 V_hig
+ 6.361010000e-07 V_hig
+ 6.362000000e-07 V_hig
+ 6.362010000e-07 V_hig
+ 6.363000000e-07 V_hig
+ 6.363010000e-07 V_hig
+ 6.364000000e-07 V_hig
+ 6.364010000e-07 V_hig
+ 6.365000000e-07 V_hig
+ 6.365010000e-07 V_hig
+ 6.366000000e-07 V_hig
+ 6.366010000e-07 V_hig
+ 6.367000000e-07 V_hig
+ 6.367010000e-07 V_hig
+ 6.368000000e-07 V_hig
+ 6.368010000e-07 V_hig
+ 6.369000000e-07 V_hig
+ 6.369010000e-07 V_low
+ 6.370000000e-07 V_low
+ 6.370010000e-07 V_low
+ 6.371000000e-07 V_low
+ 6.371010000e-07 V_low
+ 6.372000000e-07 V_low
+ 6.372010000e-07 V_low
+ 6.373000000e-07 V_low
+ 6.373010000e-07 V_low
+ 6.374000000e-07 V_low
+ 6.374010000e-07 V_low
+ 6.375000000e-07 V_low
+ 6.375010000e-07 V_low
+ 6.376000000e-07 V_low
+ 6.376010000e-07 V_low
+ 6.377000000e-07 V_low
+ 6.377010000e-07 V_low
+ 6.378000000e-07 V_low
+ 6.378010000e-07 V_low
+ 6.379000000e-07 V_low
+ 6.379010000e-07 V_low
+ 6.380000000e-07 V_low
+ 6.380010000e-07 V_low
+ 6.381000000e-07 V_low
+ 6.381010000e-07 V_low
+ 6.382000000e-07 V_low
+ 6.382010000e-07 V_low
+ 6.383000000e-07 V_low
+ 6.383010000e-07 V_low
+ 6.384000000e-07 V_low
+ 6.384010000e-07 V_low
+ 6.385000000e-07 V_low
+ 6.385010000e-07 V_low
+ 6.386000000e-07 V_low
+ 6.386010000e-07 V_low
+ 6.387000000e-07 V_low
+ 6.387010000e-07 V_low
+ 6.388000000e-07 V_low
+ 6.388010000e-07 V_low
+ 6.389000000e-07 V_low
+ 6.389010000e-07 V_low
+ 6.390000000e-07 V_low
+ 6.390010000e-07 V_low
+ 6.391000000e-07 V_low
+ 6.391010000e-07 V_low
+ 6.392000000e-07 V_low
+ 6.392010000e-07 V_low
+ 6.393000000e-07 V_low
+ 6.393010000e-07 V_low
+ 6.394000000e-07 V_low
+ 6.394010000e-07 V_low
+ 6.395000000e-07 V_low
+ 6.395010000e-07 V_low
+ 6.396000000e-07 V_low
+ 6.396010000e-07 V_low
+ 6.397000000e-07 V_low
+ 6.397010000e-07 V_low
+ 6.398000000e-07 V_low
+ 6.398010000e-07 V_low
+ 6.399000000e-07 V_low
+ 6.399010000e-07 V_low
+ 6.400000000e-07 V_low
+ 6.400010000e-07 V_low
+ 6.401000000e-07 V_low
+ 6.401010000e-07 V_low
+ 6.402000000e-07 V_low
+ 6.402010000e-07 V_low
+ 6.403000000e-07 V_low
+ 6.403010000e-07 V_low
+ 6.404000000e-07 V_low
+ 6.404010000e-07 V_low
+ 6.405000000e-07 V_low
+ 6.405010000e-07 V_low
+ 6.406000000e-07 V_low
+ 6.406010000e-07 V_low
+ 6.407000000e-07 V_low
+ 6.407010000e-07 V_low
+ 6.408000000e-07 V_low
+ 6.408010000e-07 V_low
+ 6.409000000e-07 V_low
+ 6.409010000e-07 V_hig
+ 6.410000000e-07 V_hig
+ 6.410010000e-07 V_hig
+ 6.411000000e-07 V_hig
+ 6.411010000e-07 V_hig
+ 6.412000000e-07 V_hig
+ 6.412010000e-07 V_hig
+ 6.413000000e-07 V_hig
+ 6.413010000e-07 V_hig
+ 6.414000000e-07 V_hig
+ 6.414010000e-07 V_hig
+ 6.415000000e-07 V_hig
+ 6.415010000e-07 V_hig
+ 6.416000000e-07 V_hig
+ 6.416010000e-07 V_hig
+ 6.417000000e-07 V_hig
+ 6.417010000e-07 V_hig
+ 6.418000000e-07 V_hig
+ 6.418010000e-07 V_hig
+ 6.419000000e-07 V_hig
+ 6.419010000e-07 V_hig
+ 6.420000000e-07 V_hig
+ 6.420010000e-07 V_hig
+ 6.421000000e-07 V_hig
+ 6.421010000e-07 V_hig
+ 6.422000000e-07 V_hig
+ 6.422010000e-07 V_hig
+ 6.423000000e-07 V_hig
+ 6.423010000e-07 V_hig
+ 6.424000000e-07 V_hig
+ 6.424010000e-07 V_hig
+ 6.425000000e-07 V_hig
+ 6.425010000e-07 V_hig
+ 6.426000000e-07 V_hig
+ 6.426010000e-07 V_hig
+ 6.427000000e-07 V_hig
+ 6.427010000e-07 V_hig
+ 6.428000000e-07 V_hig
+ 6.428010000e-07 V_hig
+ 6.429000000e-07 V_hig
+ 6.429010000e-07 V_hig
+ 6.430000000e-07 V_hig
+ 6.430010000e-07 V_hig
+ 6.431000000e-07 V_hig
+ 6.431010000e-07 V_hig
+ 6.432000000e-07 V_hig
+ 6.432010000e-07 V_hig
+ 6.433000000e-07 V_hig
+ 6.433010000e-07 V_hig
+ 6.434000000e-07 V_hig
+ 6.434010000e-07 V_hig
+ 6.435000000e-07 V_hig
+ 6.435010000e-07 V_hig
+ 6.436000000e-07 V_hig
+ 6.436010000e-07 V_hig
+ 6.437000000e-07 V_hig
+ 6.437010000e-07 V_hig
+ 6.438000000e-07 V_hig
+ 6.438010000e-07 V_hig
+ 6.439000000e-07 V_hig
+ 6.439010000e-07 V_low
+ 6.440000000e-07 V_low
+ 6.440010000e-07 V_low
+ 6.441000000e-07 V_low
+ 6.441010000e-07 V_low
+ 6.442000000e-07 V_low
+ 6.442010000e-07 V_low
+ 6.443000000e-07 V_low
+ 6.443010000e-07 V_low
+ 6.444000000e-07 V_low
+ 6.444010000e-07 V_low
+ 6.445000000e-07 V_low
+ 6.445010000e-07 V_low
+ 6.446000000e-07 V_low
+ 6.446010000e-07 V_low
+ 6.447000000e-07 V_low
+ 6.447010000e-07 V_low
+ 6.448000000e-07 V_low
+ 6.448010000e-07 V_low
+ 6.449000000e-07 V_low
+ 6.449010000e-07 V_hig
+ 6.450000000e-07 V_hig
+ 6.450010000e-07 V_hig
+ 6.451000000e-07 V_hig
+ 6.451010000e-07 V_hig
+ 6.452000000e-07 V_hig
+ 6.452010000e-07 V_hig
+ 6.453000000e-07 V_hig
+ 6.453010000e-07 V_hig
+ 6.454000000e-07 V_hig
+ 6.454010000e-07 V_hig
+ 6.455000000e-07 V_hig
+ 6.455010000e-07 V_hig
+ 6.456000000e-07 V_hig
+ 6.456010000e-07 V_hig
+ 6.457000000e-07 V_hig
+ 6.457010000e-07 V_hig
+ 6.458000000e-07 V_hig
+ 6.458010000e-07 V_hig
+ 6.459000000e-07 V_hig
+ 6.459010000e-07 V_hig
+ 6.460000000e-07 V_hig
+ 6.460010000e-07 V_hig
+ 6.461000000e-07 V_hig
+ 6.461010000e-07 V_hig
+ 6.462000000e-07 V_hig
+ 6.462010000e-07 V_hig
+ 6.463000000e-07 V_hig
+ 6.463010000e-07 V_hig
+ 6.464000000e-07 V_hig
+ 6.464010000e-07 V_hig
+ 6.465000000e-07 V_hig
+ 6.465010000e-07 V_hig
+ 6.466000000e-07 V_hig
+ 6.466010000e-07 V_hig
+ 6.467000000e-07 V_hig
+ 6.467010000e-07 V_hig
+ 6.468000000e-07 V_hig
+ 6.468010000e-07 V_hig
+ 6.469000000e-07 V_hig
+ 6.469010000e-07 V_hig
+ 6.470000000e-07 V_hig
+ 6.470010000e-07 V_hig
+ 6.471000000e-07 V_hig
+ 6.471010000e-07 V_hig
+ 6.472000000e-07 V_hig
+ 6.472010000e-07 V_hig
+ 6.473000000e-07 V_hig
+ 6.473010000e-07 V_hig
+ 6.474000000e-07 V_hig
+ 6.474010000e-07 V_hig
+ 6.475000000e-07 V_hig
+ 6.475010000e-07 V_hig
+ 6.476000000e-07 V_hig
+ 6.476010000e-07 V_hig
+ 6.477000000e-07 V_hig
+ 6.477010000e-07 V_hig
+ 6.478000000e-07 V_hig
+ 6.478010000e-07 V_hig
+ 6.479000000e-07 V_hig
+ 6.479010000e-07 V_hig
+ 6.480000000e-07 V_hig
+ 6.480010000e-07 V_hig
+ 6.481000000e-07 V_hig
+ 6.481010000e-07 V_hig
+ 6.482000000e-07 V_hig
+ 6.482010000e-07 V_hig
+ 6.483000000e-07 V_hig
+ 6.483010000e-07 V_hig
+ 6.484000000e-07 V_hig
+ 6.484010000e-07 V_hig
+ 6.485000000e-07 V_hig
+ 6.485010000e-07 V_hig
+ 6.486000000e-07 V_hig
+ 6.486010000e-07 V_hig
+ 6.487000000e-07 V_hig
+ 6.487010000e-07 V_hig
+ 6.488000000e-07 V_hig
+ 6.488010000e-07 V_hig
+ 6.489000000e-07 V_hig
+ 6.489010000e-07 V_hig
+ 6.490000000e-07 V_hig
+ 6.490010000e-07 V_hig
+ 6.491000000e-07 V_hig
+ 6.491010000e-07 V_hig
+ 6.492000000e-07 V_hig
+ 6.492010000e-07 V_hig
+ 6.493000000e-07 V_hig
+ 6.493010000e-07 V_hig
+ 6.494000000e-07 V_hig
+ 6.494010000e-07 V_hig
+ 6.495000000e-07 V_hig
+ 6.495010000e-07 V_hig
+ 6.496000000e-07 V_hig
+ 6.496010000e-07 V_hig
+ 6.497000000e-07 V_hig
+ 6.497010000e-07 V_hig
+ 6.498000000e-07 V_hig
+ 6.498010000e-07 V_hig
+ 6.499000000e-07 V_hig
+ 6.499010000e-07 V_low
+ 6.500000000e-07 V_low
+ 6.500010000e-07 V_low
+ 6.501000000e-07 V_low
+ 6.501010000e-07 V_low
+ 6.502000000e-07 V_low
+ 6.502010000e-07 V_low
+ 6.503000000e-07 V_low
+ 6.503010000e-07 V_low
+ 6.504000000e-07 V_low
+ 6.504010000e-07 V_low
+ 6.505000000e-07 V_low
+ 6.505010000e-07 V_low
+ 6.506000000e-07 V_low
+ 6.506010000e-07 V_low
+ 6.507000000e-07 V_low
+ 6.507010000e-07 V_low
+ 6.508000000e-07 V_low
+ 6.508010000e-07 V_low
+ 6.509000000e-07 V_low
+ 6.509010000e-07 V_hig
+ 6.510000000e-07 V_hig
+ 6.510010000e-07 V_hig
+ 6.511000000e-07 V_hig
+ 6.511010000e-07 V_hig
+ 6.512000000e-07 V_hig
+ 6.512010000e-07 V_hig
+ 6.513000000e-07 V_hig
+ 6.513010000e-07 V_hig
+ 6.514000000e-07 V_hig
+ 6.514010000e-07 V_hig
+ 6.515000000e-07 V_hig
+ 6.515010000e-07 V_hig
+ 6.516000000e-07 V_hig
+ 6.516010000e-07 V_hig
+ 6.517000000e-07 V_hig
+ 6.517010000e-07 V_hig
+ 6.518000000e-07 V_hig
+ 6.518010000e-07 V_hig
+ 6.519000000e-07 V_hig
+ 6.519010000e-07 V_low
+ 6.520000000e-07 V_low
+ 6.520010000e-07 V_low
+ 6.521000000e-07 V_low
+ 6.521010000e-07 V_low
+ 6.522000000e-07 V_low
+ 6.522010000e-07 V_low
+ 6.523000000e-07 V_low
+ 6.523010000e-07 V_low
+ 6.524000000e-07 V_low
+ 6.524010000e-07 V_low
+ 6.525000000e-07 V_low
+ 6.525010000e-07 V_low
+ 6.526000000e-07 V_low
+ 6.526010000e-07 V_low
+ 6.527000000e-07 V_low
+ 6.527010000e-07 V_low
+ 6.528000000e-07 V_low
+ 6.528010000e-07 V_low
+ 6.529000000e-07 V_low
+ 6.529010000e-07 V_hig
+ 6.530000000e-07 V_hig
+ 6.530010000e-07 V_hig
+ 6.531000000e-07 V_hig
+ 6.531010000e-07 V_hig
+ 6.532000000e-07 V_hig
+ 6.532010000e-07 V_hig
+ 6.533000000e-07 V_hig
+ 6.533010000e-07 V_hig
+ 6.534000000e-07 V_hig
+ 6.534010000e-07 V_hig
+ 6.535000000e-07 V_hig
+ 6.535010000e-07 V_hig
+ 6.536000000e-07 V_hig
+ 6.536010000e-07 V_hig
+ 6.537000000e-07 V_hig
+ 6.537010000e-07 V_hig
+ 6.538000000e-07 V_hig
+ 6.538010000e-07 V_hig
+ 6.539000000e-07 V_hig
+ 6.539010000e-07 V_low
+ 6.540000000e-07 V_low
+ 6.540010000e-07 V_low
+ 6.541000000e-07 V_low
+ 6.541010000e-07 V_low
+ 6.542000000e-07 V_low
+ 6.542010000e-07 V_low
+ 6.543000000e-07 V_low
+ 6.543010000e-07 V_low
+ 6.544000000e-07 V_low
+ 6.544010000e-07 V_low
+ 6.545000000e-07 V_low
+ 6.545010000e-07 V_low
+ 6.546000000e-07 V_low
+ 6.546010000e-07 V_low
+ 6.547000000e-07 V_low
+ 6.547010000e-07 V_low
+ 6.548000000e-07 V_low
+ 6.548010000e-07 V_low
+ 6.549000000e-07 V_low
+ 6.549010000e-07 V_low
+ 6.550000000e-07 V_low
+ 6.550010000e-07 V_low
+ 6.551000000e-07 V_low
+ 6.551010000e-07 V_low
+ 6.552000000e-07 V_low
+ 6.552010000e-07 V_low
+ 6.553000000e-07 V_low
+ 6.553010000e-07 V_low
+ 6.554000000e-07 V_low
+ 6.554010000e-07 V_low
+ 6.555000000e-07 V_low
+ 6.555010000e-07 V_low
+ 6.556000000e-07 V_low
+ 6.556010000e-07 V_low
+ 6.557000000e-07 V_low
+ 6.557010000e-07 V_low
+ 6.558000000e-07 V_low
+ 6.558010000e-07 V_low
+ 6.559000000e-07 V_low
+ 6.559010000e-07 V_hig
+ 6.560000000e-07 V_hig
+ 6.560010000e-07 V_hig
+ 6.561000000e-07 V_hig
+ 6.561010000e-07 V_hig
+ 6.562000000e-07 V_hig
+ 6.562010000e-07 V_hig
+ 6.563000000e-07 V_hig
+ 6.563010000e-07 V_hig
+ 6.564000000e-07 V_hig
+ 6.564010000e-07 V_hig
+ 6.565000000e-07 V_hig
+ 6.565010000e-07 V_hig
+ 6.566000000e-07 V_hig
+ 6.566010000e-07 V_hig
+ 6.567000000e-07 V_hig
+ 6.567010000e-07 V_hig
+ 6.568000000e-07 V_hig
+ 6.568010000e-07 V_hig
+ 6.569000000e-07 V_hig
+ 6.569010000e-07 V_hig
+ 6.570000000e-07 V_hig
+ 6.570010000e-07 V_hig
+ 6.571000000e-07 V_hig
+ 6.571010000e-07 V_hig
+ 6.572000000e-07 V_hig
+ 6.572010000e-07 V_hig
+ 6.573000000e-07 V_hig
+ 6.573010000e-07 V_hig
+ 6.574000000e-07 V_hig
+ 6.574010000e-07 V_hig
+ 6.575000000e-07 V_hig
+ 6.575010000e-07 V_hig
+ 6.576000000e-07 V_hig
+ 6.576010000e-07 V_hig
+ 6.577000000e-07 V_hig
+ 6.577010000e-07 V_hig
+ 6.578000000e-07 V_hig
+ 6.578010000e-07 V_hig
+ 6.579000000e-07 V_hig
+ 6.579010000e-07 V_hig
+ 6.580000000e-07 V_hig
+ 6.580010000e-07 V_hig
+ 6.581000000e-07 V_hig
+ 6.581010000e-07 V_hig
+ 6.582000000e-07 V_hig
+ 6.582010000e-07 V_hig
+ 6.583000000e-07 V_hig
+ 6.583010000e-07 V_hig
+ 6.584000000e-07 V_hig
+ 6.584010000e-07 V_hig
+ 6.585000000e-07 V_hig
+ 6.585010000e-07 V_hig
+ 6.586000000e-07 V_hig
+ 6.586010000e-07 V_hig
+ 6.587000000e-07 V_hig
+ 6.587010000e-07 V_hig
+ 6.588000000e-07 V_hig
+ 6.588010000e-07 V_hig
+ 6.589000000e-07 V_hig
+ 6.589010000e-07 V_hig
+ 6.590000000e-07 V_hig
+ 6.590010000e-07 V_hig
+ 6.591000000e-07 V_hig
+ 6.591010000e-07 V_hig
+ 6.592000000e-07 V_hig
+ 6.592010000e-07 V_hig
+ 6.593000000e-07 V_hig
+ 6.593010000e-07 V_hig
+ 6.594000000e-07 V_hig
+ 6.594010000e-07 V_hig
+ 6.595000000e-07 V_hig
+ 6.595010000e-07 V_hig
+ 6.596000000e-07 V_hig
+ 6.596010000e-07 V_hig
+ 6.597000000e-07 V_hig
+ 6.597010000e-07 V_hig
+ 6.598000000e-07 V_hig
+ 6.598010000e-07 V_hig
+ 6.599000000e-07 V_hig
+ 6.599010000e-07 V_hig
+ 6.600000000e-07 V_hig
+ 6.600010000e-07 V_hig
+ 6.601000000e-07 V_hig
+ 6.601010000e-07 V_hig
+ 6.602000000e-07 V_hig
+ 6.602010000e-07 V_hig
+ 6.603000000e-07 V_hig
+ 6.603010000e-07 V_hig
+ 6.604000000e-07 V_hig
+ 6.604010000e-07 V_hig
+ 6.605000000e-07 V_hig
+ 6.605010000e-07 V_hig
+ 6.606000000e-07 V_hig
+ 6.606010000e-07 V_hig
+ 6.607000000e-07 V_hig
+ 6.607010000e-07 V_hig
+ 6.608000000e-07 V_hig
+ 6.608010000e-07 V_hig
+ 6.609000000e-07 V_hig
+ 6.609010000e-07 V_low
+ 6.610000000e-07 V_low
+ 6.610010000e-07 V_low
+ 6.611000000e-07 V_low
+ 6.611010000e-07 V_low
+ 6.612000000e-07 V_low
+ 6.612010000e-07 V_low
+ 6.613000000e-07 V_low
+ 6.613010000e-07 V_low
+ 6.614000000e-07 V_low
+ 6.614010000e-07 V_low
+ 6.615000000e-07 V_low
+ 6.615010000e-07 V_low
+ 6.616000000e-07 V_low
+ 6.616010000e-07 V_low
+ 6.617000000e-07 V_low
+ 6.617010000e-07 V_low
+ 6.618000000e-07 V_low
+ 6.618010000e-07 V_low
+ 6.619000000e-07 V_low
+ 6.619010000e-07 V_hig
+ 6.620000000e-07 V_hig
+ 6.620010000e-07 V_hig
+ 6.621000000e-07 V_hig
+ 6.621010000e-07 V_hig
+ 6.622000000e-07 V_hig
+ 6.622010000e-07 V_hig
+ 6.623000000e-07 V_hig
+ 6.623010000e-07 V_hig
+ 6.624000000e-07 V_hig
+ 6.624010000e-07 V_hig
+ 6.625000000e-07 V_hig
+ 6.625010000e-07 V_hig
+ 6.626000000e-07 V_hig
+ 6.626010000e-07 V_hig
+ 6.627000000e-07 V_hig
+ 6.627010000e-07 V_hig
+ 6.628000000e-07 V_hig
+ 6.628010000e-07 V_hig
+ 6.629000000e-07 V_hig
+ 6.629010000e-07 V_hig
+ 6.630000000e-07 V_hig
+ 6.630010000e-07 V_hig
+ 6.631000000e-07 V_hig
+ 6.631010000e-07 V_hig
+ 6.632000000e-07 V_hig
+ 6.632010000e-07 V_hig
+ 6.633000000e-07 V_hig
+ 6.633010000e-07 V_hig
+ 6.634000000e-07 V_hig
+ 6.634010000e-07 V_hig
+ 6.635000000e-07 V_hig
+ 6.635010000e-07 V_hig
+ 6.636000000e-07 V_hig
+ 6.636010000e-07 V_hig
+ 6.637000000e-07 V_hig
+ 6.637010000e-07 V_hig
+ 6.638000000e-07 V_hig
+ 6.638010000e-07 V_hig
+ 6.639000000e-07 V_hig
+ 6.639010000e-07 V_hig
+ 6.640000000e-07 V_hig
+ 6.640010000e-07 V_hig
+ 6.641000000e-07 V_hig
+ 6.641010000e-07 V_hig
+ 6.642000000e-07 V_hig
+ 6.642010000e-07 V_hig
+ 6.643000000e-07 V_hig
+ 6.643010000e-07 V_hig
+ 6.644000000e-07 V_hig
+ 6.644010000e-07 V_hig
+ 6.645000000e-07 V_hig
+ 6.645010000e-07 V_hig
+ 6.646000000e-07 V_hig
+ 6.646010000e-07 V_hig
+ 6.647000000e-07 V_hig
+ 6.647010000e-07 V_hig
+ 6.648000000e-07 V_hig
+ 6.648010000e-07 V_hig
+ 6.649000000e-07 V_hig
+ 6.649010000e-07 V_low
+ 6.650000000e-07 V_low
+ 6.650010000e-07 V_low
+ 6.651000000e-07 V_low
+ 6.651010000e-07 V_low
+ 6.652000000e-07 V_low
+ 6.652010000e-07 V_low
+ 6.653000000e-07 V_low
+ 6.653010000e-07 V_low
+ 6.654000000e-07 V_low
+ 6.654010000e-07 V_low
+ 6.655000000e-07 V_low
+ 6.655010000e-07 V_low
+ 6.656000000e-07 V_low
+ 6.656010000e-07 V_low
+ 6.657000000e-07 V_low
+ 6.657010000e-07 V_low
+ 6.658000000e-07 V_low
+ 6.658010000e-07 V_low
+ 6.659000000e-07 V_low
+ 6.659010000e-07 V_low
+ 6.660000000e-07 V_low
+ 6.660010000e-07 V_low
+ 6.661000000e-07 V_low
+ 6.661010000e-07 V_low
+ 6.662000000e-07 V_low
+ 6.662010000e-07 V_low
+ 6.663000000e-07 V_low
+ 6.663010000e-07 V_low
+ 6.664000000e-07 V_low
+ 6.664010000e-07 V_low
+ 6.665000000e-07 V_low
+ 6.665010000e-07 V_low
+ 6.666000000e-07 V_low
+ 6.666010000e-07 V_low
+ 6.667000000e-07 V_low
+ 6.667010000e-07 V_low
+ 6.668000000e-07 V_low
+ 6.668010000e-07 V_low
+ 6.669000000e-07 V_low
+ 6.669010000e-07 V_hig
+ 6.670000000e-07 V_hig
+ 6.670010000e-07 V_hig
+ 6.671000000e-07 V_hig
+ 6.671010000e-07 V_hig
+ 6.672000000e-07 V_hig
+ 6.672010000e-07 V_hig
+ 6.673000000e-07 V_hig
+ 6.673010000e-07 V_hig
+ 6.674000000e-07 V_hig
+ 6.674010000e-07 V_hig
+ 6.675000000e-07 V_hig
+ 6.675010000e-07 V_hig
+ 6.676000000e-07 V_hig
+ 6.676010000e-07 V_hig
+ 6.677000000e-07 V_hig
+ 6.677010000e-07 V_hig
+ 6.678000000e-07 V_hig
+ 6.678010000e-07 V_hig
+ 6.679000000e-07 V_hig
+ 6.679010000e-07 V_hig
+ 6.680000000e-07 V_hig
+ 6.680010000e-07 V_hig
+ 6.681000000e-07 V_hig
+ 6.681010000e-07 V_hig
+ 6.682000000e-07 V_hig
+ 6.682010000e-07 V_hig
+ 6.683000000e-07 V_hig
+ 6.683010000e-07 V_hig
+ 6.684000000e-07 V_hig
+ 6.684010000e-07 V_hig
+ 6.685000000e-07 V_hig
+ 6.685010000e-07 V_hig
+ 6.686000000e-07 V_hig
+ 6.686010000e-07 V_hig
+ 6.687000000e-07 V_hig
+ 6.687010000e-07 V_hig
+ 6.688000000e-07 V_hig
+ 6.688010000e-07 V_hig
+ 6.689000000e-07 V_hig
+ 6.689010000e-07 V_hig
+ 6.690000000e-07 V_hig
+ 6.690010000e-07 V_hig
+ 6.691000000e-07 V_hig
+ 6.691010000e-07 V_hig
+ 6.692000000e-07 V_hig
+ 6.692010000e-07 V_hig
+ 6.693000000e-07 V_hig
+ 6.693010000e-07 V_hig
+ 6.694000000e-07 V_hig
+ 6.694010000e-07 V_hig
+ 6.695000000e-07 V_hig
+ 6.695010000e-07 V_hig
+ 6.696000000e-07 V_hig
+ 6.696010000e-07 V_hig
+ 6.697000000e-07 V_hig
+ 6.697010000e-07 V_hig
+ 6.698000000e-07 V_hig
+ 6.698010000e-07 V_hig
+ 6.699000000e-07 V_hig
+ 6.699010000e-07 V_low
+ 6.700000000e-07 V_low
+ 6.700010000e-07 V_low
+ 6.701000000e-07 V_low
+ 6.701010000e-07 V_low
+ 6.702000000e-07 V_low
+ 6.702010000e-07 V_low
+ 6.703000000e-07 V_low
+ 6.703010000e-07 V_low
+ 6.704000000e-07 V_low
+ 6.704010000e-07 V_low
+ 6.705000000e-07 V_low
+ 6.705010000e-07 V_low
+ 6.706000000e-07 V_low
+ 6.706010000e-07 V_low
+ 6.707000000e-07 V_low
+ 6.707010000e-07 V_low
+ 6.708000000e-07 V_low
+ 6.708010000e-07 V_low
+ 6.709000000e-07 V_low
+ 6.709010000e-07 V_low
+ 6.710000000e-07 V_low
+ 6.710010000e-07 V_low
+ 6.711000000e-07 V_low
+ 6.711010000e-07 V_low
+ 6.712000000e-07 V_low
+ 6.712010000e-07 V_low
+ 6.713000000e-07 V_low
+ 6.713010000e-07 V_low
+ 6.714000000e-07 V_low
+ 6.714010000e-07 V_low
+ 6.715000000e-07 V_low
+ 6.715010000e-07 V_low
+ 6.716000000e-07 V_low
+ 6.716010000e-07 V_low
+ 6.717000000e-07 V_low
+ 6.717010000e-07 V_low
+ 6.718000000e-07 V_low
+ 6.718010000e-07 V_low
+ 6.719000000e-07 V_low
+ 6.719010000e-07 V_low
+ 6.720000000e-07 V_low
+ 6.720010000e-07 V_low
+ 6.721000000e-07 V_low
+ 6.721010000e-07 V_low
+ 6.722000000e-07 V_low
+ 6.722010000e-07 V_low
+ 6.723000000e-07 V_low
+ 6.723010000e-07 V_low
+ 6.724000000e-07 V_low
+ 6.724010000e-07 V_low
+ 6.725000000e-07 V_low
+ 6.725010000e-07 V_low
+ 6.726000000e-07 V_low
+ 6.726010000e-07 V_low
+ 6.727000000e-07 V_low
+ 6.727010000e-07 V_low
+ 6.728000000e-07 V_low
+ 6.728010000e-07 V_low
+ 6.729000000e-07 V_low
+ 6.729010000e-07 V_hig
+ 6.730000000e-07 V_hig
+ 6.730010000e-07 V_hig
+ 6.731000000e-07 V_hig
+ 6.731010000e-07 V_hig
+ 6.732000000e-07 V_hig
+ 6.732010000e-07 V_hig
+ 6.733000000e-07 V_hig
+ 6.733010000e-07 V_hig
+ 6.734000000e-07 V_hig
+ 6.734010000e-07 V_hig
+ 6.735000000e-07 V_hig
+ 6.735010000e-07 V_hig
+ 6.736000000e-07 V_hig
+ 6.736010000e-07 V_hig
+ 6.737000000e-07 V_hig
+ 6.737010000e-07 V_hig
+ 6.738000000e-07 V_hig
+ 6.738010000e-07 V_hig
+ 6.739000000e-07 V_hig
+ 6.739010000e-07 V_low
+ 6.740000000e-07 V_low
+ 6.740010000e-07 V_low
+ 6.741000000e-07 V_low
+ 6.741010000e-07 V_low
+ 6.742000000e-07 V_low
+ 6.742010000e-07 V_low
+ 6.743000000e-07 V_low
+ 6.743010000e-07 V_low
+ 6.744000000e-07 V_low
+ 6.744010000e-07 V_low
+ 6.745000000e-07 V_low
+ 6.745010000e-07 V_low
+ 6.746000000e-07 V_low
+ 6.746010000e-07 V_low
+ 6.747000000e-07 V_low
+ 6.747010000e-07 V_low
+ 6.748000000e-07 V_low
+ 6.748010000e-07 V_low
+ 6.749000000e-07 V_low
+ 6.749010000e-07 V_hig
+ 6.750000000e-07 V_hig
+ 6.750010000e-07 V_hig
+ 6.751000000e-07 V_hig
+ 6.751010000e-07 V_hig
+ 6.752000000e-07 V_hig
+ 6.752010000e-07 V_hig
+ 6.753000000e-07 V_hig
+ 6.753010000e-07 V_hig
+ 6.754000000e-07 V_hig
+ 6.754010000e-07 V_hig
+ 6.755000000e-07 V_hig
+ 6.755010000e-07 V_hig
+ 6.756000000e-07 V_hig
+ 6.756010000e-07 V_hig
+ 6.757000000e-07 V_hig
+ 6.757010000e-07 V_hig
+ 6.758000000e-07 V_hig
+ 6.758010000e-07 V_hig
+ 6.759000000e-07 V_hig
+ 6.759010000e-07 V_hig
+ 6.760000000e-07 V_hig
+ 6.760010000e-07 V_hig
+ 6.761000000e-07 V_hig
+ 6.761010000e-07 V_hig
+ 6.762000000e-07 V_hig
+ 6.762010000e-07 V_hig
+ 6.763000000e-07 V_hig
+ 6.763010000e-07 V_hig
+ 6.764000000e-07 V_hig
+ 6.764010000e-07 V_hig
+ 6.765000000e-07 V_hig
+ 6.765010000e-07 V_hig
+ 6.766000000e-07 V_hig
+ 6.766010000e-07 V_hig
+ 6.767000000e-07 V_hig
+ 6.767010000e-07 V_hig
+ 6.768000000e-07 V_hig
+ 6.768010000e-07 V_hig
+ 6.769000000e-07 V_hig
+ 6.769010000e-07 V_hig
+ 6.770000000e-07 V_hig
+ 6.770010000e-07 V_hig
+ 6.771000000e-07 V_hig
+ 6.771010000e-07 V_hig
+ 6.772000000e-07 V_hig
+ 6.772010000e-07 V_hig
+ 6.773000000e-07 V_hig
+ 6.773010000e-07 V_hig
+ 6.774000000e-07 V_hig
+ 6.774010000e-07 V_hig
+ 6.775000000e-07 V_hig
+ 6.775010000e-07 V_hig
+ 6.776000000e-07 V_hig
+ 6.776010000e-07 V_hig
+ 6.777000000e-07 V_hig
+ 6.777010000e-07 V_hig
+ 6.778000000e-07 V_hig
+ 6.778010000e-07 V_hig
+ 6.779000000e-07 V_hig
+ 6.779010000e-07 V_hig
+ 6.780000000e-07 V_hig
+ 6.780010000e-07 V_hig
+ 6.781000000e-07 V_hig
+ 6.781010000e-07 V_hig
+ 6.782000000e-07 V_hig
+ 6.782010000e-07 V_hig
+ 6.783000000e-07 V_hig
+ 6.783010000e-07 V_hig
+ 6.784000000e-07 V_hig
+ 6.784010000e-07 V_hig
+ 6.785000000e-07 V_hig
+ 6.785010000e-07 V_hig
+ 6.786000000e-07 V_hig
+ 6.786010000e-07 V_hig
+ 6.787000000e-07 V_hig
+ 6.787010000e-07 V_hig
+ 6.788000000e-07 V_hig
+ 6.788010000e-07 V_hig
+ 6.789000000e-07 V_hig
+ 6.789010000e-07 V_low
+ 6.790000000e-07 V_low
+ 6.790010000e-07 V_low
+ 6.791000000e-07 V_low
+ 6.791010000e-07 V_low
+ 6.792000000e-07 V_low
+ 6.792010000e-07 V_low
+ 6.793000000e-07 V_low
+ 6.793010000e-07 V_low
+ 6.794000000e-07 V_low
+ 6.794010000e-07 V_low
+ 6.795000000e-07 V_low
+ 6.795010000e-07 V_low
+ 6.796000000e-07 V_low
+ 6.796010000e-07 V_low
+ 6.797000000e-07 V_low
+ 6.797010000e-07 V_low
+ 6.798000000e-07 V_low
+ 6.798010000e-07 V_low
+ 6.799000000e-07 V_low
+ 6.799010000e-07 V_hig
+ 6.800000000e-07 V_hig
+ 6.800010000e-07 V_hig
+ 6.801000000e-07 V_hig
+ 6.801010000e-07 V_hig
+ 6.802000000e-07 V_hig
+ 6.802010000e-07 V_hig
+ 6.803000000e-07 V_hig
+ 6.803010000e-07 V_hig
+ 6.804000000e-07 V_hig
+ 6.804010000e-07 V_hig
+ 6.805000000e-07 V_hig
+ 6.805010000e-07 V_hig
+ 6.806000000e-07 V_hig
+ 6.806010000e-07 V_hig
+ 6.807000000e-07 V_hig
+ 6.807010000e-07 V_hig
+ 6.808000000e-07 V_hig
+ 6.808010000e-07 V_hig
+ 6.809000000e-07 V_hig
+ 6.809010000e-07 V_low
+ 6.810000000e-07 V_low
+ 6.810010000e-07 V_low
+ 6.811000000e-07 V_low
+ 6.811010000e-07 V_low
+ 6.812000000e-07 V_low
+ 6.812010000e-07 V_low
+ 6.813000000e-07 V_low
+ 6.813010000e-07 V_low
+ 6.814000000e-07 V_low
+ 6.814010000e-07 V_low
+ 6.815000000e-07 V_low
+ 6.815010000e-07 V_low
+ 6.816000000e-07 V_low
+ 6.816010000e-07 V_low
+ 6.817000000e-07 V_low
+ 6.817010000e-07 V_low
+ 6.818000000e-07 V_low
+ 6.818010000e-07 V_low
+ 6.819000000e-07 V_low
+ 6.819010000e-07 V_low
+ 6.820000000e-07 V_low
+ 6.820010000e-07 V_low
+ 6.821000000e-07 V_low
+ 6.821010000e-07 V_low
+ 6.822000000e-07 V_low
+ 6.822010000e-07 V_low
+ 6.823000000e-07 V_low
+ 6.823010000e-07 V_low
+ 6.824000000e-07 V_low
+ 6.824010000e-07 V_low
+ 6.825000000e-07 V_low
+ 6.825010000e-07 V_low
+ 6.826000000e-07 V_low
+ 6.826010000e-07 V_low
+ 6.827000000e-07 V_low
+ 6.827010000e-07 V_low
+ 6.828000000e-07 V_low
+ 6.828010000e-07 V_low
+ 6.829000000e-07 V_low
+ 6.829010000e-07 V_hig
+ 6.830000000e-07 V_hig
+ 6.830010000e-07 V_hig
+ 6.831000000e-07 V_hig
+ 6.831010000e-07 V_hig
+ 6.832000000e-07 V_hig
+ 6.832010000e-07 V_hig
+ 6.833000000e-07 V_hig
+ 6.833010000e-07 V_hig
+ 6.834000000e-07 V_hig
+ 6.834010000e-07 V_hig
+ 6.835000000e-07 V_hig
+ 6.835010000e-07 V_hig
+ 6.836000000e-07 V_hig
+ 6.836010000e-07 V_hig
+ 6.837000000e-07 V_hig
+ 6.837010000e-07 V_hig
+ 6.838000000e-07 V_hig
+ 6.838010000e-07 V_hig
+ 6.839000000e-07 V_hig
+ 6.839010000e-07 V_hig
+ 6.840000000e-07 V_hig
+ 6.840010000e-07 V_hig
+ 6.841000000e-07 V_hig
+ 6.841010000e-07 V_hig
+ 6.842000000e-07 V_hig
+ 6.842010000e-07 V_hig
+ 6.843000000e-07 V_hig
+ 6.843010000e-07 V_hig
+ 6.844000000e-07 V_hig
+ 6.844010000e-07 V_hig
+ 6.845000000e-07 V_hig
+ 6.845010000e-07 V_hig
+ 6.846000000e-07 V_hig
+ 6.846010000e-07 V_hig
+ 6.847000000e-07 V_hig
+ 6.847010000e-07 V_hig
+ 6.848000000e-07 V_hig
+ 6.848010000e-07 V_hig
+ 6.849000000e-07 V_hig
+ 6.849010000e-07 V_hig
+ 6.850000000e-07 V_hig
+ 6.850010000e-07 V_hig
+ 6.851000000e-07 V_hig
+ 6.851010000e-07 V_hig
+ 6.852000000e-07 V_hig
+ 6.852010000e-07 V_hig
+ 6.853000000e-07 V_hig
+ 6.853010000e-07 V_hig
+ 6.854000000e-07 V_hig
+ 6.854010000e-07 V_hig
+ 6.855000000e-07 V_hig
+ 6.855010000e-07 V_hig
+ 6.856000000e-07 V_hig
+ 6.856010000e-07 V_hig
+ 6.857000000e-07 V_hig
+ 6.857010000e-07 V_hig
+ 6.858000000e-07 V_hig
+ 6.858010000e-07 V_hig
+ 6.859000000e-07 V_hig
+ 6.859010000e-07 V_low
+ 6.860000000e-07 V_low
+ 6.860010000e-07 V_low
+ 6.861000000e-07 V_low
+ 6.861010000e-07 V_low
+ 6.862000000e-07 V_low
+ 6.862010000e-07 V_low
+ 6.863000000e-07 V_low
+ 6.863010000e-07 V_low
+ 6.864000000e-07 V_low
+ 6.864010000e-07 V_low
+ 6.865000000e-07 V_low
+ 6.865010000e-07 V_low
+ 6.866000000e-07 V_low
+ 6.866010000e-07 V_low
+ 6.867000000e-07 V_low
+ 6.867010000e-07 V_low
+ 6.868000000e-07 V_low
+ 6.868010000e-07 V_low
+ 6.869000000e-07 V_low
+ 6.869010000e-07 V_hig
+ 6.870000000e-07 V_hig
+ 6.870010000e-07 V_hig
+ 6.871000000e-07 V_hig
+ 6.871010000e-07 V_hig
+ 6.872000000e-07 V_hig
+ 6.872010000e-07 V_hig
+ 6.873000000e-07 V_hig
+ 6.873010000e-07 V_hig
+ 6.874000000e-07 V_hig
+ 6.874010000e-07 V_hig
+ 6.875000000e-07 V_hig
+ 6.875010000e-07 V_hig
+ 6.876000000e-07 V_hig
+ 6.876010000e-07 V_hig
+ 6.877000000e-07 V_hig
+ 6.877010000e-07 V_hig
+ 6.878000000e-07 V_hig
+ 6.878010000e-07 V_hig
+ 6.879000000e-07 V_hig
+ 6.879010000e-07 V_hig
+ 6.880000000e-07 V_hig
+ 6.880010000e-07 V_hig
+ 6.881000000e-07 V_hig
+ 6.881010000e-07 V_hig
+ 6.882000000e-07 V_hig
+ 6.882010000e-07 V_hig
+ 6.883000000e-07 V_hig
+ 6.883010000e-07 V_hig
+ 6.884000000e-07 V_hig
+ 6.884010000e-07 V_hig
+ 6.885000000e-07 V_hig
+ 6.885010000e-07 V_hig
+ 6.886000000e-07 V_hig
+ 6.886010000e-07 V_hig
+ 6.887000000e-07 V_hig
+ 6.887010000e-07 V_hig
+ 6.888000000e-07 V_hig
+ 6.888010000e-07 V_hig
+ 6.889000000e-07 V_hig
+ 6.889010000e-07 V_low
+ 6.890000000e-07 V_low
+ 6.890010000e-07 V_low
+ 6.891000000e-07 V_low
+ 6.891010000e-07 V_low
+ 6.892000000e-07 V_low
+ 6.892010000e-07 V_low
+ 6.893000000e-07 V_low
+ 6.893010000e-07 V_low
+ 6.894000000e-07 V_low
+ 6.894010000e-07 V_low
+ 6.895000000e-07 V_low
+ 6.895010000e-07 V_low
+ 6.896000000e-07 V_low
+ 6.896010000e-07 V_low
+ 6.897000000e-07 V_low
+ 6.897010000e-07 V_low
+ 6.898000000e-07 V_low
+ 6.898010000e-07 V_low
+ 6.899000000e-07 V_low
+ 6.899010000e-07 V_low
+ 6.900000000e-07 V_low
+ 6.900010000e-07 V_low
+ 6.901000000e-07 V_low
+ 6.901010000e-07 V_low
+ 6.902000000e-07 V_low
+ 6.902010000e-07 V_low
+ 6.903000000e-07 V_low
+ 6.903010000e-07 V_low
+ 6.904000000e-07 V_low
+ 6.904010000e-07 V_low
+ 6.905000000e-07 V_low
+ 6.905010000e-07 V_low
+ 6.906000000e-07 V_low
+ 6.906010000e-07 V_low
+ 6.907000000e-07 V_low
+ 6.907010000e-07 V_low
+ 6.908000000e-07 V_low
+ 6.908010000e-07 V_low
+ 6.909000000e-07 V_low
+ 6.909010000e-07 V_low
+ 6.910000000e-07 V_low
+ 6.910010000e-07 V_low
+ 6.911000000e-07 V_low
+ 6.911010000e-07 V_low
+ 6.912000000e-07 V_low
+ 6.912010000e-07 V_low
+ 6.913000000e-07 V_low
+ 6.913010000e-07 V_low
+ 6.914000000e-07 V_low
+ 6.914010000e-07 V_low
+ 6.915000000e-07 V_low
+ 6.915010000e-07 V_low
+ 6.916000000e-07 V_low
+ 6.916010000e-07 V_low
+ 6.917000000e-07 V_low
+ 6.917010000e-07 V_low
+ 6.918000000e-07 V_low
+ 6.918010000e-07 V_low
+ 6.919000000e-07 V_low
+ 6.919010000e-07 V_low
+ 6.920000000e-07 V_low
+ 6.920010000e-07 V_low
+ 6.921000000e-07 V_low
+ 6.921010000e-07 V_low
+ 6.922000000e-07 V_low
+ 6.922010000e-07 V_low
+ 6.923000000e-07 V_low
+ 6.923010000e-07 V_low
+ 6.924000000e-07 V_low
+ 6.924010000e-07 V_low
+ 6.925000000e-07 V_low
+ 6.925010000e-07 V_low
+ 6.926000000e-07 V_low
+ 6.926010000e-07 V_low
+ 6.927000000e-07 V_low
+ 6.927010000e-07 V_low
+ 6.928000000e-07 V_low
+ 6.928010000e-07 V_low
+ 6.929000000e-07 V_low
+ 6.929010000e-07 V_low
+ 6.930000000e-07 V_low
+ 6.930010000e-07 V_low
+ 6.931000000e-07 V_low
+ 6.931010000e-07 V_low
+ 6.932000000e-07 V_low
+ 6.932010000e-07 V_low
+ 6.933000000e-07 V_low
+ 6.933010000e-07 V_low
+ 6.934000000e-07 V_low
+ 6.934010000e-07 V_low
+ 6.935000000e-07 V_low
+ 6.935010000e-07 V_low
+ 6.936000000e-07 V_low
+ 6.936010000e-07 V_low
+ 6.937000000e-07 V_low
+ 6.937010000e-07 V_low
+ 6.938000000e-07 V_low
+ 6.938010000e-07 V_low
+ 6.939000000e-07 V_low
+ 6.939010000e-07 V_low
+ 6.940000000e-07 V_low
+ 6.940010000e-07 V_low
+ 6.941000000e-07 V_low
+ 6.941010000e-07 V_low
+ 6.942000000e-07 V_low
+ 6.942010000e-07 V_low
+ 6.943000000e-07 V_low
+ 6.943010000e-07 V_low
+ 6.944000000e-07 V_low
+ 6.944010000e-07 V_low
+ 6.945000000e-07 V_low
+ 6.945010000e-07 V_low
+ 6.946000000e-07 V_low
+ 6.946010000e-07 V_low
+ 6.947000000e-07 V_low
+ 6.947010000e-07 V_low
+ 6.948000000e-07 V_low
+ 6.948010000e-07 V_low
+ 6.949000000e-07 V_low
+ 6.949010000e-07 V_low
+ 6.950000000e-07 V_low
+ 6.950010000e-07 V_low
+ 6.951000000e-07 V_low
+ 6.951010000e-07 V_low
+ 6.952000000e-07 V_low
+ 6.952010000e-07 V_low
+ 6.953000000e-07 V_low
+ 6.953010000e-07 V_low
+ 6.954000000e-07 V_low
+ 6.954010000e-07 V_low
+ 6.955000000e-07 V_low
+ 6.955010000e-07 V_low
+ 6.956000000e-07 V_low
+ 6.956010000e-07 V_low
+ 6.957000000e-07 V_low
+ 6.957010000e-07 V_low
+ 6.958000000e-07 V_low
+ 6.958010000e-07 V_low
+ 6.959000000e-07 V_low
+ 6.959010000e-07 V_low
+ 6.960000000e-07 V_low
+ 6.960010000e-07 V_low
+ 6.961000000e-07 V_low
+ 6.961010000e-07 V_low
+ 6.962000000e-07 V_low
+ 6.962010000e-07 V_low
+ 6.963000000e-07 V_low
+ 6.963010000e-07 V_low
+ 6.964000000e-07 V_low
+ 6.964010000e-07 V_low
+ 6.965000000e-07 V_low
+ 6.965010000e-07 V_low
+ 6.966000000e-07 V_low
+ 6.966010000e-07 V_low
+ 6.967000000e-07 V_low
+ 6.967010000e-07 V_low
+ 6.968000000e-07 V_low
+ 6.968010000e-07 V_low
+ 6.969000000e-07 V_low
+ 6.969010000e-07 V_low
+ 6.970000000e-07 V_low
+ 6.970010000e-07 V_low
+ 6.971000000e-07 V_low
+ 6.971010000e-07 V_low
+ 6.972000000e-07 V_low
+ 6.972010000e-07 V_low
+ 6.973000000e-07 V_low
+ 6.973010000e-07 V_low
+ 6.974000000e-07 V_low
+ 6.974010000e-07 V_low
+ 6.975000000e-07 V_low
+ 6.975010000e-07 V_low
+ 6.976000000e-07 V_low
+ 6.976010000e-07 V_low
+ 6.977000000e-07 V_low
+ 6.977010000e-07 V_low
+ 6.978000000e-07 V_low
+ 6.978010000e-07 V_low
+ 6.979000000e-07 V_low
+ 6.979010000e-07 V_low
+ 6.980000000e-07 V_low
+ 6.980010000e-07 V_low
+ 6.981000000e-07 V_low
+ 6.981010000e-07 V_low
+ 6.982000000e-07 V_low
+ 6.982010000e-07 V_low
+ 6.983000000e-07 V_low
+ 6.983010000e-07 V_low
+ 6.984000000e-07 V_low
+ 6.984010000e-07 V_low
+ 6.985000000e-07 V_low
+ 6.985010000e-07 V_low
+ 6.986000000e-07 V_low
+ 6.986010000e-07 V_low
+ 6.987000000e-07 V_low
+ 6.987010000e-07 V_low
+ 6.988000000e-07 V_low
+ 6.988010000e-07 V_low
+ 6.989000000e-07 V_low
+ 6.989010000e-07 V_hig
+ 6.990000000e-07 V_hig
+ 6.990010000e-07 V_hig
+ 6.991000000e-07 V_hig
+ 6.991010000e-07 V_hig
+ 6.992000000e-07 V_hig
+ 6.992010000e-07 V_hig
+ 6.993000000e-07 V_hig
+ 6.993010000e-07 V_hig
+ 6.994000000e-07 V_hig
+ 6.994010000e-07 V_hig
+ 6.995000000e-07 V_hig
+ 6.995010000e-07 V_hig
+ 6.996000000e-07 V_hig
+ 6.996010000e-07 V_hig
+ 6.997000000e-07 V_hig
+ 6.997010000e-07 V_hig
+ 6.998000000e-07 V_hig
+ 6.998010000e-07 V_hig
+ 6.999000000e-07 V_hig
+ 6.999010000e-07 V_hig
+ 7.000000000e-07 V_hig
+ 7.000010000e-07 V_hig
+ 7.001000000e-07 V_hig
+ 7.001010000e-07 V_hig
+ 7.002000000e-07 V_hig
+ 7.002010000e-07 V_hig
+ 7.003000000e-07 V_hig
+ 7.003010000e-07 V_hig
+ 7.004000000e-07 V_hig
+ 7.004010000e-07 V_hig
+ 7.005000000e-07 V_hig
+ 7.005010000e-07 V_hig
+ 7.006000000e-07 V_hig
+ 7.006010000e-07 V_hig
+ 7.007000000e-07 V_hig
+ 7.007010000e-07 V_hig
+ 7.008000000e-07 V_hig
+ 7.008010000e-07 V_hig
+ 7.009000000e-07 V_hig
+ 7.009010000e-07 V_hig
+ 7.010000000e-07 V_hig
+ 7.010010000e-07 V_hig
+ 7.011000000e-07 V_hig
+ 7.011010000e-07 V_hig
+ 7.012000000e-07 V_hig
+ 7.012010000e-07 V_hig
+ 7.013000000e-07 V_hig
+ 7.013010000e-07 V_hig
+ 7.014000000e-07 V_hig
+ 7.014010000e-07 V_hig
+ 7.015000000e-07 V_hig
+ 7.015010000e-07 V_hig
+ 7.016000000e-07 V_hig
+ 7.016010000e-07 V_hig
+ 7.017000000e-07 V_hig
+ 7.017010000e-07 V_hig
+ 7.018000000e-07 V_hig
+ 7.018010000e-07 V_hig
+ 7.019000000e-07 V_hig
+ 7.019010000e-07 V_low
+ 7.020000000e-07 V_low
+ 7.020010000e-07 V_low
+ 7.021000000e-07 V_low
+ 7.021010000e-07 V_low
+ 7.022000000e-07 V_low
+ 7.022010000e-07 V_low
+ 7.023000000e-07 V_low
+ 7.023010000e-07 V_low
+ 7.024000000e-07 V_low
+ 7.024010000e-07 V_low
+ 7.025000000e-07 V_low
+ 7.025010000e-07 V_low
+ 7.026000000e-07 V_low
+ 7.026010000e-07 V_low
+ 7.027000000e-07 V_low
+ 7.027010000e-07 V_low
+ 7.028000000e-07 V_low
+ 7.028010000e-07 V_low
+ 7.029000000e-07 V_low
+ 7.029010000e-07 V_hig
+ 7.030000000e-07 V_hig
+ 7.030010000e-07 V_hig
+ 7.031000000e-07 V_hig
+ 7.031010000e-07 V_hig
+ 7.032000000e-07 V_hig
+ 7.032010000e-07 V_hig
+ 7.033000000e-07 V_hig
+ 7.033010000e-07 V_hig
+ 7.034000000e-07 V_hig
+ 7.034010000e-07 V_hig
+ 7.035000000e-07 V_hig
+ 7.035010000e-07 V_hig
+ 7.036000000e-07 V_hig
+ 7.036010000e-07 V_hig
+ 7.037000000e-07 V_hig
+ 7.037010000e-07 V_hig
+ 7.038000000e-07 V_hig
+ 7.038010000e-07 V_hig
+ 7.039000000e-07 V_hig
+ 7.039010000e-07 V_hig
+ 7.040000000e-07 V_hig
+ 7.040010000e-07 V_hig
+ 7.041000000e-07 V_hig
+ 7.041010000e-07 V_hig
+ 7.042000000e-07 V_hig
+ 7.042010000e-07 V_hig
+ 7.043000000e-07 V_hig
+ 7.043010000e-07 V_hig
+ 7.044000000e-07 V_hig
+ 7.044010000e-07 V_hig
+ 7.045000000e-07 V_hig
+ 7.045010000e-07 V_hig
+ 7.046000000e-07 V_hig
+ 7.046010000e-07 V_hig
+ 7.047000000e-07 V_hig
+ 7.047010000e-07 V_hig
+ 7.048000000e-07 V_hig
+ 7.048010000e-07 V_hig
+ 7.049000000e-07 V_hig
+ 7.049010000e-07 V_low
+ 7.050000000e-07 V_low
+ 7.050010000e-07 V_low
+ 7.051000000e-07 V_low
+ 7.051010000e-07 V_low
+ 7.052000000e-07 V_low
+ 7.052010000e-07 V_low
+ 7.053000000e-07 V_low
+ 7.053010000e-07 V_low
+ 7.054000000e-07 V_low
+ 7.054010000e-07 V_low
+ 7.055000000e-07 V_low
+ 7.055010000e-07 V_low
+ 7.056000000e-07 V_low
+ 7.056010000e-07 V_low
+ 7.057000000e-07 V_low
+ 7.057010000e-07 V_low
+ 7.058000000e-07 V_low
+ 7.058010000e-07 V_low
+ 7.059000000e-07 V_low
+ 7.059010000e-07 V_hig
+ 7.060000000e-07 V_hig
+ 7.060010000e-07 V_hig
+ 7.061000000e-07 V_hig
+ 7.061010000e-07 V_hig
+ 7.062000000e-07 V_hig
+ 7.062010000e-07 V_hig
+ 7.063000000e-07 V_hig
+ 7.063010000e-07 V_hig
+ 7.064000000e-07 V_hig
+ 7.064010000e-07 V_hig
+ 7.065000000e-07 V_hig
+ 7.065010000e-07 V_hig
+ 7.066000000e-07 V_hig
+ 7.066010000e-07 V_hig
+ 7.067000000e-07 V_hig
+ 7.067010000e-07 V_hig
+ 7.068000000e-07 V_hig
+ 7.068010000e-07 V_hig
+ 7.069000000e-07 V_hig
+ 7.069010000e-07 V_low
+ 7.070000000e-07 V_low
+ 7.070010000e-07 V_low
+ 7.071000000e-07 V_low
+ 7.071010000e-07 V_low
+ 7.072000000e-07 V_low
+ 7.072010000e-07 V_low
+ 7.073000000e-07 V_low
+ 7.073010000e-07 V_low
+ 7.074000000e-07 V_low
+ 7.074010000e-07 V_low
+ 7.075000000e-07 V_low
+ 7.075010000e-07 V_low
+ 7.076000000e-07 V_low
+ 7.076010000e-07 V_low
+ 7.077000000e-07 V_low
+ 7.077010000e-07 V_low
+ 7.078000000e-07 V_low
+ 7.078010000e-07 V_low
+ 7.079000000e-07 V_low
+ 7.079010000e-07 V_hig
+ 7.080000000e-07 V_hig
+ 7.080010000e-07 V_hig
+ 7.081000000e-07 V_hig
+ 7.081010000e-07 V_hig
+ 7.082000000e-07 V_hig
+ 7.082010000e-07 V_hig
+ 7.083000000e-07 V_hig
+ 7.083010000e-07 V_hig
+ 7.084000000e-07 V_hig
+ 7.084010000e-07 V_hig
+ 7.085000000e-07 V_hig
+ 7.085010000e-07 V_hig
+ 7.086000000e-07 V_hig
+ 7.086010000e-07 V_hig
+ 7.087000000e-07 V_hig
+ 7.087010000e-07 V_hig
+ 7.088000000e-07 V_hig
+ 7.088010000e-07 V_hig
+ 7.089000000e-07 V_hig
+ 7.089010000e-07 V_hig
+ 7.090000000e-07 V_hig
+ 7.090010000e-07 V_hig
+ 7.091000000e-07 V_hig
+ 7.091010000e-07 V_hig
+ 7.092000000e-07 V_hig
+ 7.092010000e-07 V_hig
+ 7.093000000e-07 V_hig
+ 7.093010000e-07 V_hig
+ 7.094000000e-07 V_hig
+ 7.094010000e-07 V_hig
+ 7.095000000e-07 V_hig
+ 7.095010000e-07 V_hig
+ 7.096000000e-07 V_hig
+ 7.096010000e-07 V_hig
+ 7.097000000e-07 V_hig
+ 7.097010000e-07 V_hig
+ 7.098000000e-07 V_hig
+ 7.098010000e-07 V_hig
+ 7.099000000e-07 V_hig
+ 7.099010000e-07 V_hig
+ 7.100000000e-07 V_hig
+ 7.100010000e-07 V_hig
+ 7.101000000e-07 V_hig
+ 7.101010000e-07 V_hig
+ 7.102000000e-07 V_hig
+ 7.102010000e-07 V_hig
+ 7.103000000e-07 V_hig
+ 7.103010000e-07 V_hig
+ 7.104000000e-07 V_hig
+ 7.104010000e-07 V_hig
+ 7.105000000e-07 V_hig
+ 7.105010000e-07 V_hig
+ 7.106000000e-07 V_hig
+ 7.106010000e-07 V_hig
+ 7.107000000e-07 V_hig
+ 7.107010000e-07 V_hig
+ 7.108000000e-07 V_hig
+ 7.108010000e-07 V_hig
+ 7.109000000e-07 V_hig
+ 7.109010000e-07 V_low
+ 7.110000000e-07 V_low
+ 7.110010000e-07 V_low
+ 7.111000000e-07 V_low
+ 7.111010000e-07 V_low
+ 7.112000000e-07 V_low
+ 7.112010000e-07 V_low
+ 7.113000000e-07 V_low
+ 7.113010000e-07 V_low
+ 7.114000000e-07 V_low
+ 7.114010000e-07 V_low
+ 7.115000000e-07 V_low
+ 7.115010000e-07 V_low
+ 7.116000000e-07 V_low
+ 7.116010000e-07 V_low
+ 7.117000000e-07 V_low
+ 7.117010000e-07 V_low
+ 7.118000000e-07 V_low
+ 7.118010000e-07 V_low
+ 7.119000000e-07 V_low
+ 7.119010000e-07 V_low
+ 7.120000000e-07 V_low
+ 7.120010000e-07 V_low
+ 7.121000000e-07 V_low
+ 7.121010000e-07 V_low
+ 7.122000000e-07 V_low
+ 7.122010000e-07 V_low
+ 7.123000000e-07 V_low
+ 7.123010000e-07 V_low
+ 7.124000000e-07 V_low
+ 7.124010000e-07 V_low
+ 7.125000000e-07 V_low
+ 7.125010000e-07 V_low
+ 7.126000000e-07 V_low
+ 7.126010000e-07 V_low
+ 7.127000000e-07 V_low
+ 7.127010000e-07 V_low
+ 7.128000000e-07 V_low
+ 7.128010000e-07 V_low
+ 7.129000000e-07 V_low
+ 7.129010000e-07 V_low
+ 7.130000000e-07 V_low
+ 7.130010000e-07 V_low
+ 7.131000000e-07 V_low
+ 7.131010000e-07 V_low
+ 7.132000000e-07 V_low
+ 7.132010000e-07 V_low
+ 7.133000000e-07 V_low
+ 7.133010000e-07 V_low
+ 7.134000000e-07 V_low
+ 7.134010000e-07 V_low
+ 7.135000000e-07 V_low
+ 7.135010000e-07 V_low
+ 7.136000000e-07 V_low
+ 7.136010000e-07 V_low
+ 7.137000000e-07 V_low
+ 7.137010000e-07 V_low
+ 7.138000000e-07 V_low
+ 7.138010000e-07 V_low
+ 7.139000000e-07 V_low
+ 7.139010000e-07 V_low
+ 7.140000000e-07 V_low
+ 7.140010000e-07 V_low
+ 7.141000000e-07 V_low
+ 7.141010000e-07 V_low
+ 7.142000000e-07 V_low
+ 7.142010000e-07 V_low
+ 7.143000000e-07 V_low
+ 7.143010000e-07 V_low
+ 7.144000000e-07 V_low
+ 7.144010000e-07 V_low
+ 7.145000000e-07 V_low
+ 7.145010000e-07 V_low
+ 7.146000000e-07 V_low
+ 7.146010000e-07 V_low
+ 7.147000000e-07 V_low
+ 7.147010000e-07 V_low
+ 7.148000000e-07 V_low
+ 7.148010000e-07 V_low
+ 7.149000000e-07 V_low
+ 7.149010000e-07 V_low
+ 7.150000000e-07 V_low
+ 7.150010000e-07 V_low
+ 7.151000000e-07 V_low
+ 7.151010000e-07 V_low
+ 7.152000000e-07 V_low
+ 7.152010000e-07 V_low
+ 7.153000000e-07 V_low
+ 7.153010000e-07 V_low
+ 7.154000000e-07 V_low
+ 7.154010000e-07 V_low
+ 7.155000000e-07 V_low
+ 7.155010000e-07 V_low
+ 7.156000000e-07 V_low
+ 7.156010000e-07 V_low
+ 7.157000000e-07 V_low
+ 7.157010000e-07 V_low
+ 7.158000000e-07 V_low
+ 7.158010000e-07 V_low
+ 7.159000000e-07 V_low
+ 7.159010000e-07 V_hig
+ 7.160000000e-07 V_hig
+ 7.160010000e-07 V_hig
+ 7.161000000e-07 V_hig
+ 7.161010000e-07 V_hig
+ 7.162000000e-07 V_hig
+ 7.162010000e-07 V_hig
+ 7.163000000e-07 V_hig
+ 7.163010000e-07 V_hig
+ 7.164000000e-07 V_hig
+ 7.164010000e-07 V_hig
+ 7.165000000e-07 V_hig
+ 7.165010000e-07 V_hig
+ 7.166000000e-07 V_hig
+ 7.166010000e-07 V_hig
+ 7.167000000e-07 V_hig
+ 7.167010000e-07 V_hig
+ 7.168000000e-07 V_hig
+ 7.168010000e-07 V_hig
+ 7.169000000e-07 V_hig
+ 7.169010000e-07 V_low
+ 7.170000000e-07 V_low
+ 7.170010000e-07 V_low
+ 7.171000000e-07 V_low
+ 7.171010000e-07 V_low
+ 7.172000000e-07 V_low
+ 7.172010000e-07 V_low
+ 7.173000000e-07 V_low
+ 7.173010000e-07 V_low
+ 7.174000000e-07 V_low
+ 7.174010000e-07 V_low
+ 7.175000000e-07 V_low
+ 7.175010000e-07 V_low
+ 7.176000000e-07 V_low
+ 7.176010000e-07 V_low
+ 7.177000000e-07 V_low
+ 7.177010000e-07 V_low
+ 7.178000000e-07 V_low
+ 7.178010000e-07 V_low
+ 7.179000000e-07 V_low
+ 7.179010000e-07 V_low
+ 7.180000000e-07 V_low
+ 7.180010000e-07 V_low
+ 7.181000000e-07 V_low
+ 7.181010000e-07 V_low
+ 7.182000000e-07 V_low
+ 7.182010000e-07 V_low
+ 7.183000000e-07 V_low
+ 7.183010000e-07 V_low
+ 7.184000000e-07 V_low
+ 7.184010000e-07 V_low
+ 7.185000000e-07 V_low
+ 7.185010000e-07 V_low
+ 7.186000000e-07 V_low
+ 7.186010000e-07 V_low
+ 7.187000000e-07 V_low
+ 7.187010000e-07 V_low
+ 7.188000000e-07 V_low
+ 7.188010000e-07 V_low
+ 7.189000000e-07 V_low
+ 7.189010000e-07 V_low
+ 7.190000000e-07 V_low
+ 7.190010000e-07 V_low
+ 7.191000000e-07 V_low
+ 7.191010000e-07 V_low
+ 7.192000000e-07 V_low
+ 7.192010000e-07 V_low
+ 7.193000000e-07 V_low
+ 7.193010000e-07 V_low
+ 7.194000000e-07 V_low
+ 7.194010000e-07 V_low
+ 7.195000000e-07 V_low
+ 7.195010000e-07 V_low
+ 7.196000000e-07 V_low
+ 7.196010000e-07 V_low
+ 7.197000000e-07 V_low
+ 7.197010000e-07 V_low
+ 7.198000000e-07 V_low
+ 7.198010000e-07 V_low
+ 7.199000000e-07 V_low
+ 7.199010000e-07 V_hig
+ 7.200000000e-07 V_hig
+ 7.200010000e-07 V_hig
+ 7.201000000e-07 V_hig
+ 7.201010000e-07 V_hig
+ 7.202000000e-07 V_hig
+ 7.202010000e-07 V_hig
+ 7.203000000e-07 V_hig
+ 7.203010000e-07 V_hig
+ 7.204000000e-07 V_hig
+ 7.204010000e-07 V_hig
+ 7.205000000e-07 V_hig
+ 7.205010000e-07 V_hig
+ 7.206000000e-07 V_hig
+ 7.206010000e-07 V_hig
+ 7.207000000e-07 V_hig
+ 7.207010000e-07 V_hig
+ 7.208000000e-07 V_hig
+ 7.208010000e-07 V_hig
+ 7.209000000e-07 V_hig
+ 7.209010000e-07 V_low
+ 7.210000000e-07 V_low
+ 7.210010000e-07 V_low
+ 7.211000000e-07 V_low
+ 7.211010000e-07 V_low
+ 7.212000000e-07 V_low
+ 7.212010000e-07 V_low
+ 7.213000000e-07 V_low
+ 7.213010000e-07 V_low
+ 7.214000000e-07 V_low
+ 7.214010000e-07 V_low
+ 7.215000000e-07 V_low
+ 7.215010000e-07 V_low
+ 7.216000000e-07 V_low
+ 7.216010000e-07 V_low
+ 7.217000000e-07 V_low
+ 7.217010000e-07 V_low
+ 7.218000000e-07 V_low
+ 7.218010000e-07 V_low
+ 7.219000000e-07 V_low
+ 7.219010000e-07 V_low
+ 7.220000000e-07 V_low
+ 7.220010000e-07 V_low
+ 7.221000000e-07 V_low
+ 7.221010000e-07 V_low
+ 7.222000000e-07 V_low
+ 7.222010000e-07 V_low
+ 7.223000000e-07 V_low
+ 7.223010000e-07 V_low
+ 7.224000000e-07 V_low
+ 7.224010000e-07 V_low
+ 7.225000000e-07 V_low
+ 7.225010000e-07 V_low
+ 7.226000000e-07 V_low
+ 7.226010000e-07 V_low
+ 7.227000000e-07 V_low
+ 7.227010000e-07 V_low
+ 7.228000000e-07 V_low
+ 7.228010000e-07 V_low
+ 7.229000000e-07 V_low
+ 7.229010000e-07 V_low
+ 7.230000000e-07 V_low
+ 7.230010000e-07 V_low
+ 7.231000000e-07 V_low
+ 7.231010000e-07 V_low
+ 7.232000000e-07 V_low
+ 7.232010000e-07 V_low
+ 7.233000000e-07 V_low
+ 7.233010000e-07 V_low
+ 7.234000000e-07 V_low
+ 7.234010000e-07 V_low
+ 7.235000000e-07 V_low
+ 7.235010000e-07 V_low
+ 7.236000000e-07 V_low
+ 7.236010000e-07 V_low
+ 7.237000000e-07 V_low
+ 7.237010000e-07 V_low
+ 7.238000000e-07 V_low
+ 7.238010000e-07 V_low
+ 7.239000000e-07 V_low
+ 7.239010000e-07 V_low
+ 7.240000000e-07 V_low
+ 7.240010000e-07 V_low
+ 7.241000000e-07 V_low
+ 7.241010000e-07 V_low
+ 7.242000000e-07 V_low
+ 7.242010000e-07 V_low
+ 7.243000000e-07 V_low
+ 7.243010000e-07 V_low
+ 7.244000000e-07 V_low
+ 7.244010000e-07 V_low
+ 7.245000000e-07 V_low
+ 7.245010000e-07 V_low
+ 7.246000000e-07 V_low
+ 7.246010000e-07 V_low
+ 7.247000000e-07 V_low
+ 7.247010000e-07 V_low
+ 7.248000000e-07 V_low
+ 7.248010000e-07 V_low
+ 7.249000000e-07 V_low
+ 7.249010000e-07 V_low
+ 7.250000000e-07 V_low
+ 7.250010000e-07 V_low
+ 7.251000000e-07 V_low
+ 7.251010000e-07 V_low
+ 7.252000000e-07 V_low
+ 7.252010000e-07 V_low
+ 7.253000000e-07 V_low
+ 7.253010000e-07 V_low
+ 7.254000000e-07 V_low
+ 7.254010000e-07 V_low
+ 7.255000000e-07 V_low
+ 7.255010000e-07 V_low
+ 7.256000000e-07 V_low
+ 7.256010000e-07 V_low
+ 7.257000000e-07 V_low
+ 7.257010000e-07 V_low
+ 7.258000000e-07 V_low
+ 7.258010000e-07 V_low
+ 7.259000000e-07 V_low
+ 7.259010000e-07 V_hig
+ 7.260000000e-07 V_hig
+ 7.260010000e-07 V_hig
+ 7.261000000e-07 V_hig
+ 7.261010000e-07 V_hig
+ 7.262000000e-07 V_hig
+ 7.262010000e-07 V_hig
+ 7.263000000e-07 V_hig
+ 7.263010000e-07 V_hig
+ 7.264000000e-07 V_hig
+ 7.264010000e-07 V_hig
+ 7.265000000e-07 V_hig
+ 7.265010000e-07 V_hig
+ 7.266000000e-07 V_hig
+ 7.266010000e-07 V_hig
+ 7.267000000e-07 V_hig
+ 7.267010000e-07 V_hig
+ 7.268000000e-07 V_hig
+ 7.268010000e-07 V_hig
+ 7.269000000e-07 V_hig
+ 7.269010000e-07 V_hig
+ 7.270000000e-07 V_hig
+ 7.270010000e-07 V_hig
+ 7.271000000e-07 V_hig
+ 7.271010000e-07 V_hig
+ 7.272000000e-07 V_hig
+ 7.272010000e-07 V_hig
+ 7.273000000e-07 V_hig
+ 7.273010000e-07 V_hig
+ 7.274000000e-07 V_hig
+ 7.274010000e-07 V_hig
+ 7.275000000e-07 V_hig
+ 7.275010000e-07 V_hig
+ 7.276000000e-07 V_hig
+ 7.276010000e-07 V_hig
+ 7.277000000e-07 V_hig
+ 7.277010000e-07 V_hig
+ 7.278000000e-07 V_hig
+ 7.278010000e-07 V_hig
+ 7.279000000e-07 V_hig
+ 7.279010000e-07 V_low
+ 7.280000000e-07 V_low
+ 7.280010000e-07 V_low
+ 7.281000000e-07 V_low
+ 7.281010000e-07 V_low
+ 7.282000000e-07 V_low
+ 7.282010000e-07 V_low
+ 7.283000000e-07 V_low
+ 7.283010000e-07 V_low
+ 7.284000000e-07 V_low
+ 7.284010000e-07 V_low
+ 7.285000000e-07 V_low
+ 7.285010000e-07 V_low
+ 7.286000000e-07 V_low
+ 7.286010000e-07 V_low
+ 7.287000000e-07 V_low
+ 7.287010000e-07 V_low
+ 7.288000000e-07 V_low
+ 7.288010000e-07 V_low
+ 7.289000000e-07 V_low
+ 7.289010000e-07 V_hig
+ 7.290000000e-07 V_hig
+ 7.290010000e-07 V_hig
+ 7.291000000e-07 V_hig
+ 7.291010000e-07 V_hig
+ 7.292000000e-07 V_hig
+ 7.292010000e-07 V_hig
+ 7.293000000e-07 V_hig
+ 7.293010000e-07 V_hig
+ 7.294000000e-07 V_hig
+ 7.294010000e-07 V_hig
+ 7.295000000e-07 V_hig
+ 7.295010000e-07 V_hig
+ 7.296000000e-07 V_hig
+ 7.296010000e-07 V_hig
+ 7.297000000e-07 V_hig
+ 7.297010000e-07 V_hig
+ 7.298000000e-07 V_hig
+ 7.298010000e-07 V_hig
+ 7.299000000e-07 V_hig
+ 7.299010000e-07 V_low
+ 7.300000000e-07 V_low
+ 7.300010000e-07 V_low
+ 7.301000000e-07 V_low
+ 7.301010000e-07 V_low
+ 7.302000000e-07 V_low
+ 7.302010000e-07 V_low
+ 7.303000000e-07 V_low
+ 7.303010000e-07 V_low
+ 7.304000000e-07 V_low
+ 7.304010000e-07 V_low
+ 7.305000000e-07 V_low
+ 7.305010000e-07 V_low
+ 7.306000000e-07 V_low
+ 7.306010000e-07 V_low
+ 7.307000000e-07 V_low
+ 7.307010000e-07 V_low
+ 7.308000000e-07 V_low
+ 7.308010000e-07 V_low
+ 7.309000000e-07 V_low
+ 7.309010000e-07 V_hig
+ 7.310000000e-07 V_hig
+ 7.310010000e-07 V_hig
+ 7.311000000e-07 V_hig
+ 7.311010000e-07 V_hig
+ 7.312000000e-07 V_hig
+ 7.312010000e-07 V_hig
+ 7.313000000e-07 V_hig
+ 7.313010000e-07 V_hig
+ 7.314000000e-07 V_hig
+ 7.314010000e-07 V_hig
+ 7.315000000e-07 V_hig
+ 7.315010000e-07 V_hig
+ 7.316000000e-07 V_hig
+ 7.316010000e-07 V_hig
+ 7.317000000e-07 V_hig
+ 7.317010000e-07 V_hig
+ 7.318000000e-07 V_hig
+ 7.318010000e-07 V_hig
+ 7.319000000e-07 V_hig
+ 7.319010000e-07 V_hig
+ 7.320000000e-07 V_hig
+ 7.320010000e-07 V_hig
+ 7.321000000e-07 V_hig
+ 7.321010000e-07 V_hig
+ 7.322000000e-07 V_hig
+ 7.322010000e-07 V_hig
+ 7.323000000e-07 V_hig
+ 7.323010000e-07 V_hig
+ 7.324000000e-07 V_hig
+ 7.324010000e-07 V_hig
+ 7.325000000e-07 V_hig
+ 7.325010000e-07 V_hig
+ 7.326000000e-07 V_hig
+ 7.326010000e-07 V_hig
+ 7.327000000e-07 V_hig
+ 7.327010000e-07 V_hig
+ 7.328000000e-07 V_hig
+ 7.328010000e-07 V_hig
+ 7.329000000e-07 V_hig
+ 7.329010000e-07 V_low
+ 7.330000000e-07 V_low
+ 7.330010000e-07 V_low
+ 7.331000000e-07 V_low
+ 7.331010000e-07 V_low
+ 7.332000000e-07 V_low
+ 7.332010000e-07 V_low
+ 7.333000000e-07 V_low
+ 7.333010000e-07 V_low
+ 7.334000000e-07 V_low
+ 7.334010000e-07 V_low
+ 7.335000000e-07 V_low
+ 7.335010000e-07 V_low
+ 7.336000000e-07 V_low
+ 7.336010000e-07 V_low
+ 7.337000000e-07 V_low
+ 7.337010000e-07 V_low
+ 7.338000000e-07 V_low
+ 7.338010000e-07 V_low
+ 7.339000000e-07 V_low
+ 7.339010000e-07 V_low
+ 7.340000000e-07 V_low
+ 7.340010000e-07 V_low
+ 7.341000000e-07 V_low
+ 7.341010000e-07 V_low
+ 7.342000000e-07 V_low
+ 7.342010000e-07 V_low
+ 7.343000000e-07 V_low
+ 7.343010000e-07 V_low
+ 7.344000000e-07 V_low
+ 7.344010000e-07 V_low
+ 7.345000000e-07 V_low
+ 7.345010000e-07 V_low
+ 7.346000000e-07 V_low
+ 7.346010000e-07 V_low
+ 7.347000000e-07 V_low
+ 7.347010000e-07 V_low
+ 7.348000000e-07 V_low
+ 7.348010000e-07 V_low
+ 7.349000000e-07 V_low
+ 7.349010000e-07 V_hig
+ 7.350000000e-07 V_hig
+ 7.350010000e-07 V_hig
+ 7.351000000e-07 V_hig
+ 7.351010000e-07 V_hig
+ 7.352000000e-07 V_hig
+ 7.352010000e-07 V_hig
+ 7.353000000e-07 V_hig
+ 7.353010000e-07 V_hig
+ 7.354000000e-07 V_hig
+ 7.354010000e-07 V_hig
+ 7.355000000e-07 V_hig
+ 7.355010000e-07 V_hig
+ 7.356000000e-07 V_hig
+ 7.356010000e-07 V_hig
+ 7.357000000e-07 V_hig
+ 7.357010000e-07 V_hig
+ 7.358000000e-07 V_hig
+ 7.358010000e-07 V_hig
+ 7.359000000e-07 V_hig
+ 7.359010000e-07 V_hig
+ 7.360000000e-07 V_hig
+ 7.360010000e-07 V_hig
+ 7.361000000e-07 V_hig
+ 7.361010000e-07 V_hig
+ 7.362000000e-07 V_hig
+ 7.362010000e-07 V_hig
+ 7.363000000e-07 V_hig
+ 7.363010000e-07 V_hig
+ 7.364000000e-07 V_hig
+ 7.364010000e-07 V_hig
+ 7.365000000e-07 V_hig
+ 7.365010000e-07 V_hig
+ 7.366000000e-07 V_hig
+ 7.366010000e-07 V_hig
+ 7.367000000e-07 V_hig
+ 7.367010000e-07 V_hig
+ 7.368000000e-07 V_hig
+ 7.368010000e-07 V_hig
+ 7.369000000e-07 V_hig
+ 7.369010000e-07 V_low
+ 7.370000000e-07 V_low
+ 7.370010000e-07 V_low
+ 7.371000000e-07 V_low
+ 7.371010000e-07 V_low
+ 7.372000000e-07 V_low
+ 7.372010000e-07 V_low
+ 7.373000000e-07 V_low
+ 7.373010000e-07 V_low
+ 7.374000000e-07 V_low
+ 7.374010000e-07 V_low
+ 7.375000000e-07 V_low
+ 7.375010000e-07 V_low
+ 7.376000000e-07 V_low
+ 7.376010000e-07 V_low
+ 7.377000000e-07 V_low
+ 7.377010000e-07 V_low
+ 7.378000000e-07 V_low
+ 7.378010000e-07 V_low
+ 7.379000000e-07 V_low
+ 7.379010000e-07 V_hig
+ 7.380000000e-07 V_hig
+ 7.380010000e-07 V_hig
+ 7.381000000e-07 V_hig
+ 7.381010000e-07 V_hig
+ 7.382000000e-07 V_hig
+ 7.382010000e-07 V_hig
+ 7.383000000e-07 V_hig
+ 7.383010000e-07 V_hig
+ 7.384000000e-07 V_hig
+ 7.384010000e-07 V_hig
+ 7.385000000e-07 V_hig
+ 7.385010000e-07 V_hig
+ 7.386000000e-07 V_hig
+ 7.386010000e-07 V_hig
+ 7.387000000e-07 V_hig
+ 7.387010000e-07 V_hig
+ 7.388000000e-07 V_hig
+ 7.388010000e-07 V_hig
+ 7.389000000e-07 V_hig
+ 7.389010000e-07 V_low
+ 7.390000000e-07 V_low
+ 7.390010000e-07 V_low
+ 7.391000000e-07 V_low
+ 7.391010000e-07 V_low
+ 7.392000000e-07 V_low
+ 7.392010000e-07 V_low
+ 7.393000000e-07 V_low
+ 7.393010000e-07 V_low
+ 7.394000000e-07 V_low
+ 7.394010000e-07 V_low
+ 7.395000000e-07 V_low
+ 7.395010000e-07 V_low
+ 7.396000000e-07 V_low
+ 7.396010000e-07 V_low
+ 7.397000000e-07 V_low
+ 7.397010000e-07 V_low
+ 7.398000000e-07 V_low
+ 7.398010000e-07 V_low
+ 7.399000000e-07 V_low
+ 7.399010000e-07 V_low
+ 7.400000000e-07 V_low
+ 7.400010000e-07 V_low
+ 7.401000000e-07 V_low
+ 7.401010000e-07 V_low
+ 7.402000000e-07 V_low
+ 7.402010000e-07 V_low
+ 7.403000000e-07 V_low
+ 7.403010000e-07 V_low
+ 7.404000000e-07 V_low
+ 7.404010000e-07 V_low
+ 7.405000000e-07 V_low
+ 7.405010000e-07 V_low
+ 7.406000000e-07 V_low
+ 7.406010000e-07 V_low
+ 7.407000000e-07 V_low
+ 7.407010000e-07 V_low
+ 7.408000000e-07 V_low
+ 7.408010000e-07 V_low
+ 7.409000000e-07 V_low
+ 7.409010000e-07 V_low
+ 7.410000000e-07 V_low
+ 7.410010000e-07 V_low
+ 7.411000000e-07 V_low
+ 7.411010000e-07 V_low
+ 7.412000000e-07 V_low
+ 7.412010000e-07 V_low
+ 7.413000000e-07 V_low
+ 7.413010000e-07 V_low
+ 7.414000000e-07 V_low
+ 7.414010000e-07 V_low
+ 7.415000000e-07 V_low
+ 7.415010000e-07 V_low
+ 7.416000000e-07 V_low
+ 7.416010000e-07 V_low
+ 7.417000000e-07 V_low
+ 7.417010000e-07 V_low
+ 7.418000000e-07 V_low
+ 7.418010000e-07 V_low
+ 7.419000000e-07 V_low
+ 7.419010000e-07 V_hig
+ 7.420000000e-07 V_hig
+ 7.420010000e-07 V_hig
+ 7.421000000e-07 V_hig
+ 7.421010000e-07 V_hig
+ 7.422000000e-07 V_hig
+ 7.422010000e-07 V_hig
+ 7.423000000e-07 V_hig
+ 7.423010000e-07 V_hig
+ 7.424000000e-07 V_hig
+ 7.424010000e-07 V_hig
+ 7.425000000e-07 V_hig
+ 7.425010000e-07 V_hig
+ 7.426000000e-07 V_hig
+ 7.426010000e-07 V_hig
+ 7.427000000e-07 V_hig
+ 7.427010000e-07 V_hig
+ 7.428000000e-07 V_hig
+ 7.428010000e-07 V_hig
+ 7.429000000e-07 V_hig
+ 7.429010000e-07 V_hig
+ 7.430000000e-07 V_hig
+ 7.430010000e-07 V_hig
+ 7.431000000e-07 V_hig
+ 7.431010000e-07 V_hig
+ 7.432000000e-07 V_hig
+ 7.432010000e-07 V_hig
+ 7.433000000e-07 V_hig
+ 7.433010000e-07 V_hig
+ 7.434000000e-07 V_hig
+ 7.434010000e-07 V_hig
+ 7.435000000e-07 V_hig
+ 7.435010000e-07 V_hig
+ 7.436000000e-07 V_hig
+ 7.436010000e-07 V_hig
+ 7.437000000e-07 V_hig
+ 7.437010000e-07 V_hig
+ 7.438000000e-07 V_hig
+ 7.438010000e-07 V_hig
+ 7.439000000e-07 V_hig
+ 7.439010000e-07 V_low
+ 7.440000000e-07 V_low
+ 7.440010000e-07 V_low
+ 7.441000000e-07 V_low
+ 7.441010000e-07 V_low
+ 7.442000000e-07 V_low
+ 7.442010000e-07 V_low
+ 7.443000000e-07 V_low
+ 7.443010000e-07 V_low
+ 7.444000000e-07 V_low
+ 7.444010000e-07 V_low
+ 7.445000000e-07 V_low
+ 7.445010000e-07 V_low
+ 7.446000000e-07 V_low
+ 7.446010000e-07 V_low
+ 7.447000000e-07 V_low
+ 7.447010000e-07 V_low
+ 7.448000000e-07 V_low
+ 7.448010000e-07 V_low
+ 7.449000000e-07 V_low
+ 7.449010000e-07 V_low
+ 7.450000000e-07 V_low
+ 7.450010000e-07 V_low
+ 7.451000000e-07 V_low
+ 7.451010000e-07 V_low
+ 7.452000000e-07 V_low
+ 7.452010000e-07 V_low
+ 7.453000000e-07 V_low
+ 7.453010000e-07 V_low
+ 7.454000000e-07 V_low
+ 7.454010000e-07 V_low
+ 7.455000000e-07 V_low
+ 7.455010000e-07 V_low
+ 7.456000000e-07 V_low
+ 7.456010000e-07 V_low
+ 7.457000000e-07 V_low
+ 7.457010000e-07 V_low
+ 7.458000000e-07 V_low
+ 7.458010000e-07 V_low
+ 7.459000000e-07 V_low
+ 7.459010000e-07 V_low
+ 7.460000000e-07 V_low
+ 7.460010000e-07 V_low
+ 7.461000000e-07 V_low
+ 7.461010000e-07 V_low
+ 7.462000000e-07 V_low
+ 7.462010000e-07 V_low
+ 7.463000000e-07 V_low
+ 7.463010000e-07 V_low
+ 7.464000000e-07 V_low
+ 7.464010000e-07 V_low
+ 7.465000000e-07 V_low
+ 7.465010000e-07 V_low
+ 7.466000000e-07 V_low
+ 7.466010000e-07 V_low
+ 7.467000000e-07 V_low
+ 7.467010000e-07 V_low
+ 7.468000000e-07 V_low
+ 7.468010000e-07 V_low
+ 7.469000000e-07 V_low
+ 7.469010000e-07 V_hig
+ 7.470000000e-07 V_hig
+ 7.470010000e-07 V_hig
+ 7.471000000e-07 V_hig
+ 7.471010000e-07 V_hig
+ 7.472000000e-07 V_hig
+ 7.472010000e-07 V_hig
+ 7.473000000e-07 V_hig
+ 7.473010000e-07 V_hig
+ 7.474000000e-07 V_hig
+ 7.474010000e-07 V_hig
+ 7.475000000e-07 V_hig
+ 7.475010000e-07 V_hig
+ 7.476000000e-07 V_hig
+ 7.476010000e-07 V_hig
+ 7.477000000e-07 V_hig
+ 7.477010000e-07 V_hig
+ 7.478000000e-07 V_hig
+ 7.478010000e-07 V_hig
+ 7.479000000e-07 V_hig
+ 7.479010000e-07 V_low
+ 7.480000000e-07 V_low
+ 7.480010000e-07 V_low
+ 7.481000000e-07 V_low
+ 7.481010000e-07 V_low
+ 7.482000000e-07 V_low
+ 7.482010000e-07 V_low
+ 7.483000000e-07 V_low
+ 7.483010000e-07 V_low
+ 7.484000000e-07 V_low
+ 7.484010000e-07 V_low
+ 7.485000000e-07 V_low
+ 7.485010000e-07 V_low
+ 7.486000000e-07 V_low
+ 7.486010000e-07 V_low
+ 7.487000000e-07 V_low
+ 7.487010000e-07 V_low
+ 7.488000000e-07 V_low
+ 7.488010000e-07 V_low
+ 7.489000000e-07 V_low
+ 7.489010000e-07 V_hig
+ 7.490000000e-07 V_hig
+ 7.490010000e-07 V_hig
+ 7.491000000e-07 V_hig
+ 7.491010000e-07 V_hig
+ 7.492000000e-07 V_hig
+ 7.492010000e-07 V_hig
+ 7.493000000e-07 V_hig
+ 7.493010000e-07 V_hig
+ 7.494000000e-07 V_hig
+ 7.494010000e-07 V_hig
+ 7.495000000e-07 V_hig
+ 7.495010000e-07 V_hig
+ 7.496000000e-07 V_hig
+ 7.496010000e-07 V_hig
+ 7.497000000e-07 V_hig
+ 7.497010000e-07 V_hig
+ 7.498000000e-07 V_hig
+ 7.498010000e-07 V_hig
+ 7.499000000e-07 V_hig
+ 7.499010000e-07 V_hig
+ 7.500000000e-07 V_hig
+ 7.500010000e-07 V_hig
+ 7.501000000e-07 V_hig
+ 7.501010000e-07 V_hig
+ 7.502000000e-07 V_hig
+ 7.502010000e-07 V_hig
+ 7.503000000e-07 V_hig
+ 7.503010000e-07 V_hig
+ 7.504000000e-07 V_hig
+ 7.504010000e-07 V_hig
+ 7.505000000e-07 V_hig
+ 7.505010000e-07 V_hig
+ 7.506000000e-07 V_hig
+ 7.506010000e-07 V_hig
+ 7.507000000e-07 V_hig
+ 7.507010000e-07 V_hig
+ 7.508000000e-07 V_hig
+ 7.508010000e-07 V_hig
+ 7.509000000e-07 V_hig
+ 7.509010000e-07 V_hig
+ 7.510000000e-07 V_hig
+ 7.510010000e-07 V_hig
+ 7.511000000e-07 V_hig
+ 7.511010000e-07 V_hig
+ 7.512000000e-07 V_hig
+ 7.512010000e-07 V_hig
+ 7.513000000e-07 V_hig
+ 7.513010000e-07 V_hig
+ 7.514000000e-07 V_hig
+ 7.514010000e-07 V_hig
+ 7.515000000e-07 V_hig
+ 7.515010000e-07 V_hig
+ 7.516000000e-07 V_hig
+ 7.516010000e-07 V_hig
+ 7.517000000e-07 V_hig
+ 7.517010000e-07 V_hig
+ 7.518000000e-07 V_hig
+ 7.518010000e-07 V_hig
+ 7.519000000e-07 V_hig
+ 7.519010000e-07 V_low
+ 7.520000000e-07 V_low
+ 7.520010000e-07 V_low
+ 7.521000000e-07 V_low
+ 7.521010000e-07 V_low
+ 7.522000000e-07 V_low
+ 7.522010000e-07 V_low
+ 7.523000000e-07 V_low
+ 7.523010000e-07 V_low
+ 7.524000000e-07 V_low
+ 7.524010000e-07 V_low
+ 7.525000000e-07 V_low
+ 7.525010000e-07 V_low
+ 7.526000000e-07 V_low
+ 7.526010000e-07 V_low
+ 7.527000000e-07 V_low
+ 7.527010000e-07 V_low
+ 7.528000000e-07 V_low
+ 7.528010000e-07 V_low
+ 7.529000000e-07 V_low
+ 7.529010000e-07 V_low
+ 7.530000000e-07 V_low
+ 7.530010000e-07 V_low
+ 7.531000000e-07 V_low
+ 7.531010000e-07 V_low
+ 7.532000000e-07 V_low
+ 7.532010000e-07 V_low
+ 7.533000000e-07 V_low
+ 7.533010000e-07 V_low
+ 7.534000000e-07 V_low
+ 7.534010000e-07 V_low
+ 7.535000000e-07 V_low
+ 7.535010000e-07 V_low
+ 7.536000000e-07 V_low
+ 7.536010000e-07 V_low
+ 7.537000000e-07 V_low
+ 7.537010000e-07 V_low
+ 7.538000000e-07 V_low
+ 7.538010000e-07 V_low
+ 7.539000000e-07 V_low
+ 7.539010000e-07 V_low
+ 7.540000000e-07 V_low
+ 7.540010000e-07 V_low
+ 7.541000000e-07 V_low
+ 7.541010000e-07 V_low
+ 7.542000000e-07 V_low
+ 7.542010000e-07 V_low
+ 7.543000000e-07 V_low
+ 7.543010000e-07 V_low
+ 7.544000000e-07 V_low
+ 7.544010000e-07 V_low
+ 7.545000000e-07 V_low
+ 7.545010000e-07 V_low
+ 7.546000000e-07 V_low
+ 7.546010000e-07 V_low
+ 7.547000000e-07 V_low
+ 7.547010000e-07 V_low
+ 7.548000000e-07 V_low
+ 7.548010000e-07 V_low
+ 7.549000000e-07 V_low
+ 7.549010000e-07 V_low
+ 7.550000000e-07 V_low
+ 7.550010000e-07 V_low
+ 7.551000000e-07 V_low
+ 7.551010000e-07 V_low
+ 7.552000000e-07 V_low
+ 7.552010000e-07 V_low
+ 7.553000000e-07 V_low
+ 7.553010000e-07 V_low
+ 7.554000000e-07 V_low
+ 7.554010000e-07 V_low
+ 7.555000000e-07 V_low
+ 7.555010000e-07 V_low
+ 7.556000000e-07 V_low
+ 7.556010000e-07 V_low
+ 7.557000000e-07 V_low
+ 7.557010000e-07 V_low
+ 7.558000000e-07 V_low
+ 7.558010000e-07 V_low
+ 7.559000000e-07 V_low
+ 7.559010000e-07 V_low
+ 7.560000000e-07 V_low
+ 7.560010000e-07 V_low
+ 7.561000000e-07 V_low
+ 7.561010000e-07 V_low
+ 7.562000000e-07 V_low
+ 7.562010000e-07 V_low
+ 7.563000000e-07 V_low
+ 7.563010000e-07 V_low
+ 7.564000000e-07 V_low
+ 7.564010000e-07 V_low
+ 7.565000000e-07 V_low
+ 7.565010000e-07 V_low
+ 7.566000000e-07 V_low
+ 7.566010000e-07 V_low
+ 7.567000000e-07 V_low
+ 7.567010000e-07 V_low
+ 7.568000000e-07 V_low
+ 7.568010000e-07 V_low
+ 7.569000000e-07 V_low
+ 7.569010000e-07 V_low
+ 7.570000000e-07 V_low
+ 7.570010000e-07 V_low
+ 7.571000000e-07 V_low
+ 7.571010000e-07 V_low
+ 7.572000000e-07 V_low
+ 7.572010000e-07 V_low
+ 7.573000000e-07 V_low
+ 7.573010000e-07 V_low
+ 7.574000000e-07 V_low
+ 7.574010000e-07 V_low
+ 7.575000000e-07 V_low
+ 7.575010000e-07 V_low
+ 7.576000000e-07 V_low
+ 7.576010000e-07 V_low
+ 7.577000000e-07 V_low
+ 7.577010000e-07 V_low
+ 7.578000000e-07 V_low
+ 7.578010000e-07 V_low
+ 7.579000000e-07 V_low
+ 7.579010000e-07 V_hig
+ 7.580000000e-07 V_hig
+ 7.580010000e-07 V_hig
+ 7.581000000e-07 V_hig
+ 7.581010000e-07 V_hig
+ 7.582000000e-07 V_hig
+ 7.582010000e-07 V_hig
+ 7.583000000e-07 V_hig
+ 7.583010000e-07 V_hig
+ 7.584000000e-07 V_hig
+ 7.584010000e-07 V_hig
+ 7.585000000e-07 V_hig
+ 7.585010000e-07 V_hig
+ 7.586000000e-07 V_hig
+ 7.586010000e-07 V_hig
+ 7.587000000e-07 V_hig
+ 7.587010000e-07 V_hig
+ 7.588000000e-07 V_hig
+ 7.588010000e-07 V_hig
+ 7.589000000e-07 V_hig
+ 7.589010000e-07 V_hig
+ 7.590000000e-07 V_hig
+ 7.590010000e-07 V_hig
+ 7.591000000e-07 V_hig
+ 7.591010000e-07 V_hig
+ 7.592000000e-07 V_hig
+ 7.592010000e-07 V_hig
+ 7.593000000e-07 V_hig
+ 7.593010000e-07 V_hig
+ 7.594000000e-07 V_hig
+ 7.594010000e-07 V_hig
+ 7.595000000e-07 V_hig
+ 7.595010000e-07 V_hig
+ 7.596000000e-07 V_hig
+ 7.596010000e-07 V_hig
+ 7.597000000e-07 V_hig
+ 7.597010000e-07 V_hig
+ 7.598000000e-07 V_hig
+ 7.598010000e-07 V_hig
+ 7.599000000e-07 V_hig
+ 7.599010000e-07 V_hig
+ 7.600000000e-07 V_hig
+ 7.600010000e-07 V_hig
+ 7.601000000e-07 V_hig
+ 7.601010000e-07 V_hig
+ 7.602000000e-07 V_hig
+ 7.602010000e-07 V_hig
+ 7.603000000e-07 V_hig
+ 7.603010000e-07 V_hig
+ 7.604000000e-07 V_hig
+ 7.604010000e-07 V_hig
+ 7.605000000e-07 V_hig
+ 7.605010000e-07 V_hig
+ 7.606000000e-07 V_hig
+ 7.606010000e-07 V_hig
+ 7.607000000e-07 V_hig
+ 7.607010000e-07 V_hig
+ 7.608000000e-07 V_hig
+ 7.608010000e-07 V_hig
+ 7.609000000e-07 V_hig
+ 7.609010000e-07 V_low
+ 7.610000000e-07 V_low
+ 7.610010000e-07 V_low
+ 7.611000000e-07 V_low
+ 7.611010000e-07 V_low
+ 7.612000000e-07 V_low
+ 7.612010000e-07 V_low
+ 7.613000000e-07 V_low
+ 7.613010000e-07 V_low
+ 7.614000000e-07 V_low
+ 7.614010000e-07 V_low
+ 7.615000000e-07 V_low
+ 7.615010000e-07 V_low
+ 7.616000000e-07 V_low
+ 7.616010000e-07 V_low
+ 7.617000000e-07 V_low
+ 7.617010000e-07 V_low
+ 7.618000000e-07 V_low
+ 7.618010000e-07 V_low
+ 7.619000000e-07 V_low
+ 7.619010000e-07 V_low
+ 7.620000000e-07 V_low
+ 7.620010000e-07 V_low
+ 7.621000000e-07 V_low
+ 7.621010000e-07 V_low
+ 7.622000000e-07 V_low
+ 7.622010000e-07 V_low
+ 7.623000000e-07 V_low
+ 7.623010000e-07 V_low
+ 7.624000000e-07 V_low
+ 7.624010000e-07 V_low
+ 7.625000000e-07 V_low
+ 7.625010000e-07 V_low
+ 7.626000000e-07 V_low
+ 7.626010000e-07 V_low
+ 7.627000000e-07 V_low
+ 7.627010000e-07 V_low
+ 7.628000000e-07 V_low
+ 7.628010000e-07 V_low
+ 7.629000000e-07 V_low
+ 7.629010000e-07 V_low
+ 7.630000000e-07 V_low
+ 7.630010000e-07 V_low
+ 7.631000000e-07 V_low
+ 7.631010000e-07 V_low
+ 7.632000000e-07 V_low
+ 7.632010000e-07 V_low
+ 7.633000000e-07 V_low
+ 7.633010000e-07 V_low
+ 7.634000000e-07 V_low
+ 7.634010000e-07 V_low
+ 7.635000000e-07 V_low
+ 7.635010000e-07 V_low
+ 7.636000000e-07 V_low
+ 7.636010000e-07 V_low
+ 7.637000000e-07 V_low
+ 7.637010000e-07 V_low
+ 7.638000000e-07 V_low
+ 7.638010000e-07 V_low
+ 7.639000000e-07 V_low
+ 7.639010000e-07 V_low
+ 7.640000000e-07 V_low
+ 7.640010000e-07 V_low
+ 7.641000000e-07 V_low
+ 7.641010000e-07 V_low
+ 7.642000000e-07 V_low
+ 7.642010000e-07 V_low
+ 7.643000000e-07 V_low
+ 7.643010000e-07 V_low
+ 7.644000000e-07 V_low
+ 7.644010000e-07 V_low
+ 7.645000000e-07 V_low
+ 7.645010000e-07 V_low
+ 7.646000000e-07 V_low
+ 7.646010000e-07 V_low
+ 7.647000000e-07 V_low
+ 7.647010000e-07 V_low
+ 7.648000000e-07 V_low
+ 7.648010000e-07 V_low
+ 7.649000000e-07 V_low
+ 7.649010000e-07 V_hig
+ 7.650000000e-07 V_hig
+ 7.650010000e-07 V_hig
+ 7.651000000e-07 V_hig
+ 7.651010000e-07 V_hig
+ 7.652000000e-07 V_hig
+ 7.652010000e-07 V_hig
+ 7.653000000e-07 V_hig
+ 7.653010000e-07 V_hig
+ 7.654000000e-07 V_hig
+ 7.654010000e-07 V_hig
+ 7.655000000e-07 V_hig
+ 7.655010000e-07 V_hig
+ 7.656000000e-07 V_hig
+ 7.656010000e-07 V_hig
+ 7.657000000e-07 V_hig
+ 7.657010000e-07 V_hig
+ 7.658000000e-07 V_hig
+ 7.658010000e-07 V_hig
+ 7.659000000e-07 V_hig
+ 7.659010000e-07 V_low
+ 7.660000000e-07 V_low
+ 7.660010000e-07 V_low
+ 7.661000000e-07 V_low
+ 7.661010000e-07 V_low
+ 7.662000000e-07 V_low
+ 7.662010000e-07 V_low
+ 7.663000000e-07 V_low
+ 7.663010000e-07 V_low
+ 7.664000000e-07 V_low
+ 7.664010000e-07 V_low
+ 7.665000000e-07 V_low
+ 7.665010000e-07 V_low
+ 7.666000000e-07 V_low
+ 7.666010000e-07 V_low
+ 7.667000000e-07 V_low
+ 7.667010000e-07 V_low
+ 7.668000000e-07 V_low
+ 7.668010000e-07 V_low
+ 7.669000000e-07 V_low
+ 7.669010000e-07 V_low
+ 7.670000000e-07 V_low
+ 7.670010000e-07 V_low
+ 7.671000000e-07 V_low
+ 7.671010000e-07 V_low
+ 7.672000000e-07 V_low
+ 7.672010000e-07 V_low
+ 7.673000000e-07 V_low
+ 7.673010000e-07 V_low
+ 7.674000000e-07 V_low
+ 7.674010000e-07 V_low
+ 7.675000000e-07 V_low
+ 7.675010000e-07 V_low
+ 7.676000000e-07 V_low
+ 7.676010000e-07 V_low
+ 7.677000000e-07 V_low
+ 7.677010000e-07 V_low
+ 7.678000000e-07 V_low
+ 7.678010000e-07 V_low
+ 7.679000000e-07 V_low
+ 7.679010000e-07 V_hig
+ 7.680000000e-07 V_hig
+ 7.680010000e-07 V_hig
+ 7.681000000e-07 V_hig
+ 7.681010000e-07 V_hig
+ 7.682000000e-07 V_hig
+ 7.682010000e-07 V_hig
+ 7.683000000e-07 V_hig
+ 7.683010000e-07 V_hig
+ 7.684000000e-07 V_hig
+ 7.684010000e-07 V_hig
+ 7.685000000e-07 V_hig
+ 7.685010000e-07 V_hig
+ 7.686000000e-07 V_hig
+ 7.686010000e-07 V_hig
+ 7.687000000e-07 V_hig
+ 7.687010000e-07 V_hig
+ 7.688000000e-07 V_hig
+ 7.688010000e-07 V_hig
+ 7.689000000e-07 V_hig
+ 7.689010000e-07 V_hig
+ 7.690000000e-07 V_hig
+ 7.690010000e-07 V_hig
+ 7.691000000e-07 V_hig
+ 7.691010000e-07 V_hig
+ 7.692000000e-07 V_hig
+ 7.692010000e-07 V_hig
+ 7.693000000e-07 V_hig
+ 7.693010000e-07 V_hig
+ 7.694000000e-07 V_hig
+ 7.694010000e-07 V_hig
+ 7.695000000e-07 V_hig
+ 7.695010000e-07 V_hig
+ 7.696000000e-07 V_hig
+ 7.696010000e-07 V_hig
+ 7.697000000e-07 V_hig
+ 7.697010000e-07 V_hig
+ 7.698000000e-07 V_hig
+ 7.698010000e-07 V_hig
+ 7.699000000e-07 V_hig
+ 7.699010000e-07 V_low
+ 7.700000000e-07 V_low
+ 7.700010000e-07 V_low
+ 7.701000000e-07 V_low
+ 7.701010000e-07 V_low
+ 7.702000000e-07 V_low
+ 7.702010000e-07 V_low
+ 7.703000000e-07 V_low
+ 7.703010000e-07 V_low
+ 7.704000000e-07 V_low
+ 7.704010000e-07 V_low
+ 7.705000000e-07 V_low
+ 7.705010000e-07 V_low
+ 7.706000000e-07 V_low
+ 7.706010000e-07 V_low
+ 7.707000000e-07 V_low
+ 7.707010000e-07 V_low
+ 7.708000000e-07 V_low
+ 7.708010000e-07 V_low
+ 7.709000000e-07 V_low
+ 7.709010000e-07 V_low
+ 7.710000000e-07 V_low
+ 7.710010000e-07 V_low
+ 7.711000000e-07 V_low
+ 7.711010000e-07 V_low
+ 7.712000000e-07 V_low
+ 7.712010000e-07 V_low
+ 7.713000000e-07 V_low
+ 7.713010000e-07 V_low
+ 7.714000000e-07 V_low
+ 7.714010000e-07 V_low
+ 7.715000000e-07 V_low
+ 7.715010000e-07 V_low
+ 7.716000000e-07 V_low
+ 7.716010000e-07 V_low
+ 7.717000000e-07 V_low
+ 7.717010000e-07 V_low
+ 7.718000000e-07 V_low
+ 7.718010000e-07 V_low
+ 7.719000000e-07 V_low
+ 7.719010000e-07 V_low
+ 7.720000000e-07 V_low
+ 7.720010000e-07 V_low
+ 7.721000000e-07 V_low
+ 7.721010000e-07 V_low
+ 7.722000000e-07 V_low
+ 7.722010000e-07 V_low
+ 7.723000000e-07 V_low
+ 7.723010000e-07 V_low
+ 7.724000000e-07 V_low
+ 7.724010000e-07 V_low
+ 7.725000000e-07 V_low
+ 7.725010000e-07 V_low
+ 7.726000000e-07 V_low
+ 7.726010000e-07 V_low
+ 7.727000000e-07 V_low
+ 7.727010000e-07 V_low
+ 7.728000000e-07 V_low
+ 7.728010000e-07 V_low
+ 7.729000000e-07 V_low
+ 7.729010000e-07 V_low
+ 7.730000000e-07 V_low
+ 7.730010000e-07 V_low
+ 7.731000000e-07 V_low
+ 7.731010000e-07 V_low
+ 7.732000000e-07 V_low
+ 7.732010000e-07 V_low
+ 7.733000000e-07 V_low
+ 7.733010000e-07 V_low
+ 7.734000000e-07 V_low
+ 7.734010000e-07 V_low
+ 7.735000000e-07 V_low
+ 7.735010000e-07 V_low
+ 7.736000000e-07 V_low
+ 7.736010000e-07 V_low
+ 7.737000000e-07 V_low
+ 7.737010000e-07 V_low
+ 7.738000000e-07 V_low
+ 7.738010000e-07 V_low
+ 7.739000000e-07 V_low
+ 7.739010000e-07 V_low
+ 7.740000000e-07 V_low
+ 7.740010000e-07 V_low
+ 7.741000000e-07 V_low
+ 7.741010000e-07 V_low
+ 7.742000000e-07 V_low
+ 7.742010000e-07 V_low
+ 7.743000000e-07 V_low
+ 7.743010000e-07 V_low
+ 7.744000000e-07 V_low
+ 7.744010000e-07 V_low
+ 7.745000000e-07 V_low
+ 7.745010000e-07 V_low
+ 7.746000000e-07 V_low
+ 7.746010000e-07 V_low
+ 7.747000000e-07 V_low
+ 7.747010000e-07 V_low
+ 7.748000000e-07 V_low
+ 7.748010000e-07 V_low
+ 7.749000000e-07 V_low
+ 7.749010000e-07 V_hig
+ 7.750000000e-07 V_hig
+ 7.750010000e-07 V_hig
+ 7.751000000e-07 V_hig
+ 7.751010000e-07 V_hig
+ 7.752000000e-07 V_hig
+ 7.752010000e-07 V_hig
+ 7.753000000e-07 V_hig
+ 7.753010000e-07 V_hig
+ 7.754000000e-07 V_hig
+ 7.754010000e-07 V_hig
+ 7.755000000e-07 V_hig
+ 7.755010000e-07 V_hig
+ 7.756000000e-07 V_hig
+ 7.756010000e-07 V_hig
+ 7.757000000e-07 V_hig
+ 7.757010000e-07 V_hig
+ 7.758000000e-07 V_hig
+ 7.758010000e-07 V_hig
+ 7.759000000e-07 V_hig
+ 7.759010000e-07 V_low
+ 7.760000000e-07 V_low
+ 7.760010000e-07 V_low
+ 7.761000000e-07 V_low
+ 7.761010000e-07 V_low
+ 7.762000000e-07 V_low
+ 7.762010000e-07 V_low
+ 7.763000000e-07 V_low
+ 7.763010000e-07 V_low
+ 7.764000000e-07 V_low
+ 7.764010000e-07 V_low
+ 7.765000000e-07 V_low
+ 7.765010000e-07 V_low
+ 7.766000000e-07 V_low
+ 7.766010000e-07 V_low
+ 7.767000000e-07 V_low
+ 7.767010000e-07 V_low
+ 7.768000000e-07 V_low
+ 7.768010000e-07 V_low
+ 7.769000000e-07 V_low
+ 7.769010000e-07 V_hig
+ 7.770000000e-07 V_hig
+ 7.770010000e-07 V_hig
+ 7.771000000e-07 V_hig
+ 7.771010000e-07 V_hig
+ 7.772000000e-07 V_hig
+ 7.772010000e-07 V_hig
+ 7.773000000e-07 V_hig
+ 7.773010000e-07 V_hig
+ 7.774000000e-07 V_hig
+ 7.774010000e-07 V_hig
+ 7.775000000e-07 V_hig
+ 7.775010000e-07 V_hig
+ 7.776000000e-07 V_hig
+ 7.776010000e-07 V_hig
+ 7.777000000e-07 V_hig
+ 7.777010000e-07 V_hig
+ 7.778000000e-07 V_hig
+ 7.778010000e-07 V_hig
+ 7.779000000e-07 V_hig
+ 7.779010000e-07 V_low
+ 7.780000000e-07 V_low
+ 7.780010000e-07 V_low
+ 7.781000000e-07 V_low
+ 7.781010000e-07 V_low
+ 7.782000000e-07 V_low
+ 7.782010000e-07 V_low
+ 7.783000000e-07 V_low
+ 7.783010000e-07 V_low
+ 7.784000000e-07 V_low
+ 7.784010000e-07 V_low
+ 7.785000000e-07 V_low
+ 7.785010000e-07 V_low
+ 7.786000000e-07 V_low
+ 7.786010000e-07 V_low
+ 7.787000000e-07 V_low
+ 7.787010000e-07 V_low
+ 7.788000000e-07 V_low
+ 7.788010000e-07 V_low
+ 7.789000000e-07 V_low
+ 7.789010000e-07 V_hig
+ 7.790000000e-07 V_hig
+ 7.790010000e-07 V_hig
+ 7.791000000e-07 V_hig
+ 7.791010000e-07 V_hig
+ 7.792000000e-07 V_hig
+ 7.792010000e-07 V_hig
+ 7.793000000e-07 V_hig
+ 7.793010000e-07 V_hig
+ 7.794000000e-07 V_hig
+ 7.794010000e-07 V_hig
+ 7.795000000e-07 V_hig
+ 7.795010000e-07 V_hig
+ 7.796000000e-07 V_hig
+ 7.796010000e-07 V_hig
+ 7.797000000e-07 V_hig
+ 7.797010000e-07 V_hig
+ 7.798000000e-07 V_hig
+ 7.798010000e-07 V_hig
+ 7.799000000e-07 V_hig
+ 7.799010000e-07 V_low
+ 7.800000000e-07 V_low
+ 7.800010000e-07 V_low
+ 7.801000000e-07 V_low
+ 7.801010000e-07 V_low
+ 7.802000000e-07 V_low
+ 7.802010000e-07 V_low
+ 7.803000000e-07 V_low
+ 7.803010000e-07 V_low
+ 7.804000000e-07 V_low
+ 7.804010000e-07 V_low
+ 7.805000000e-07 V_low
+ 7.805010000e-07 V_low
+ 7.806000000e-07 V_low
+ 7.806010000e-07 V_low
+ 7.807000000e-07 V_low
+ 7.807010000e-07 V_low
+ 7.808000000e-07 V_low
+ 7.808010000e-07 V_low
+ 7.809000000e-07 V_low
+ 7.809010000e-07 V_hig
+ 7.810000000e-07 V_hig
+ 7.810010000e-07 V_hig
+ 7.811000000e-07 V_hig
+ 7.811010000e-07 V_hig
+ 7.812000000e-07 V_hig
+ 7.812010000e-07 V_hig
+ 7.813000000e-07 V_hig
+ 7.813010000e-07 V_hig
+ 7.814000000e-07 V_hig
+ 7.814010000e-07 V_hig
+ 7.815000000e-07 V_hig
+ 7.815010000e-07 V_hig
+ 7.816000000e-07 V_hig
+ 7.816010000e-07 V_hig
+ 7.817000000e-07 V_hig
+ 7.817010000e-07 V_hig
+ 7.818000000e-07 V_hig
+ 7.818010000e-07 V_hig
+ 7.819000000e-07 V_hig
+ 7.819010000e-07 V_low
+ 7.820000000e-07 V_low
+ 7.820010000e-07 V_low
+ 7.821000000e-07 V_low
+ 7.821010000e-07 V_low
+ 7.822000000e-07 V_low
+ 7.822010000e-07 V_low
+ 7.823000000e-07 V_low
+ 7.823010000e-07 V_low
+ 7.824000000e-07 V_low
+ 7.824010000e-07 V_low
+ 7.825000000e-07 V_low
+ 7.825010000e-07 V_low
+ 7.826000000e-07 V_low
+ 7.826010000e-07 V_low
+ 7.827000000e-07 V_low
+ 7.827010000e-07 V_low
+ 7.828000000e-07 V_low
+ 7.828010000e-07 V_low
+ 7.829000000e-07 V_low
+ 7.829010000e-07 V_hig
+ 7.830000000e-07 V_hig
+ 7.830010000e-07 V_hig
+ 7.831000000e-07 V_hig
+ 7.831010000e-07 V_hig
+ 7.832000000e-07 V_hig
+ 7.832010000e-07 V_hig
+ 7.833000000e-07 V_hig
+ 7.833010000e-07 V_hig
+ 7.834000000e-07 V_hig
+ 7.834010000e-07 V_hig
+ 7.835000000e-07 V_hig
+ 7.835010000e-07 V_hig
+ 7.836000000e-07 V_hig
+ 7.836010000e-07 V_hig
+ 7.837000000e-07 V_hig
+ 7.837010000e-07 V_hig
+ 7.838000000e-07 V_hig
+ 7.838010000e-07 V_hig
+ 7.839000000e-07 V_hig
+ 7.839010000e-07 V_hig
+ 7.840000000e-07 V_hig
+ 7.840010000e-07 V_hig
+ 7.841000000e-07 V_hig
+ 7.841010000e-07 V_hig
+ 7.842000000e-07 V_hig
+ 7.842010000e-07 V_hig
+ 7.843000000e-07 V_hig
+ 7.843010000e-07 V_hig
+ 7.844000000e-07 V_hig
+ 7.844010000e-07 V_hig
+ 7.845000000e-07 V_hig
+ 7.845010000e-07 V_hig
+ 7.846000000e-07 V_hig
+ 7.846010000e-07 V_hig
+ 7.847000000e-07 V_hig
+ 7.847010000e-07 V_hig
+ 7.848000000e-07 V_hig
+ 7.848010000e-07 V_hig
+ 7.849000000e-07 V_hig
+ 7.849010000e-07 V_hig
+ 7.850000000e-07 V_hig
+ 7.850010000e-07 V_hig
+ 7.851000000e-07 V_hig
+ 7.851010000e-07 V_hig
+ 7.852000000e-07 V_hig
+ 7.852010000e-07 V_hig
+ 7.853000000e-07 V_hig
+ 7.853010000e-07 V_hig
+ 7.854000000e-07 V_hig
+ 7.854010000e-07 V_hig
+ 7.855000000e-07 V_hig
+ 7.855010000e-07 V_hig
+ 7.856000000e-07 V_hig
+ 7.856010000e-07 V_hig
+ 7.857000000e-07 V_hig
+ 7.857010000e-07 V_hig
+ 7.858000000e-07 V_hig
+ 7.858010000e-07 V_hig
+ 7.859000000e-07 V_hig
+ 7.859010000e-07 V_hig
+ 7.860000000e-07 V_hig
+ 7.860010000e-07 V_hig
+ 7.861000000e-07 V_hig
+ 7.861010000e-07 V_hig
+ 7.862000000e-07 V_hig
+ 7.862010000e-07 V_hig
+ 7.863000000e-07 V_hig
+ 7.863010000e-07 V_hig
+ 7.864000000e-07 V_hig
+ 7.864010000e-07 V_hig
+ 7.865000000e-07 V_hig
+ 7.865010000e-07 V_hig
+ 7.866000000e-07 V_hig
+ 7.866010000e-07 V_hig
+ 7.867000000e-07 V_hig
+ 7.867010000e-07 V_hig
+ 7.868000000e-07 V_hig
+ 7.868010000e-07 V_hig
+ 7.869000000e-07 V_hig
+ 7.869010000e-07 V_low
+ 7.870000000e-07 V_low
+ 7.870010000e-07 V_low
+ 7.871000000e-07 V_low
+ 7.871010000e-07 V_low
+ 7.872000000e-07 V_low
+ 7.872010000e-07 V_low
+ 7.873000000e-07 V_low
+ 7.873010000e-07 V_low
+ 7.874000000e-07 V_low
+ 7.874010000e-07 V_low
+ 7.875000000e-07 V_low
+ 7.875010000e-07 V_low
+ 7.876000000e-07 V_low
+ 7.876010000e-07 V_low
+ 7.877000000e-07 V_low
+ 7.877010000e-07 V_low
+ 7.878000000e-07 V_low
+ 7.878010000e-07 V_low
+ 7.879000000e-07 V_low
+ 7.879010000e-07 V_hig
+ 7.880000000e-07 V_hig
+ 7.880010000e-07 V_hig
+ 7.881000000e-07 V_hig
+ 7.881010000e-07 V_hig
+ 7.882000000e-07 V_hig
+ 7.882010000e-07 V_hig
+ 7.883000000e-07 V_hig
+ 7.883010000e-07 V_hig
+ 7.884000000e-07 V_hig
+ 7.884010000e-07 V_hig
+ 7.885000000e-07 V_hig
+ 7.885010000e-07 V_hig
+ 7.886000000e-07 V_hig
+ 7.886010000e-07 V_hig
+ 7.887000000e-07 V_hig
+ 7.887010000e-07 V_hig
+ 7.888000000e-07 V_hig
+ 7.888010000e-07 V_hig
+ 7.889000000e-07 V_hig
+ 7.889010000e-07 V_low
+ 7.890000000e-07 V_low
+ 7.890010000e-07 V_low
+ 7.891000000e-07 V_low
+ 7.891010000e-07 V_low
+ 7.892000000e-07 V_low
+ 7.892010000e-07 V_low
+ 7.893000000e-07 V_low
+ 7.893010000e-07 V_low
+ 7.894000000e-07 V_low
+ 7.894010000e-07 V_low
+ 7.895000000e-07 V_low
+ 7.895010000e-07 V_low
+ 7.896000000e-07 V_low
+ 7.896010000e-07 V_low
+ 7.897000000e-07 V_low
+ 7.897010000e-07 V_low
+ 7.898000000e-07 V_low
+ 7.898010000e-07 V_low
+ 7.899000000e-07 V_low
+ 7.899010000e-07 V_hig
+ 7.900000000e-07 V_hig
+ 7.900010000e-07 V_hig
+ 7.901000000e-07 V_hig
+ 7.901010000e-07 V_hig
+ 7.902000000e-07 V_hig
+ 7.902010000e-07 V_hig
+ 7.903000000e-07 V_hig
+ 7.903010000e-07 V_hig
+ 7.904000000e-07 V_hig
+ 7.904010000e-07 V_hig
+ 7.905000000e-07 V_hig
+ 7.905010000e-07 V_hig
+ 7.906000000e-07 V_hig
+ 7.906010000e-07 V_hig
+ 7.907000000e-07 V_hig
+ 7.907010000e-07 V_hig
+ 7.908000000e-07 V_hig
+ 7.908010000e-07 V_hig
+ 7.909000000e-07 V_hig
+ 7.909010000e-07 V_hig
+ 7.910000000e-07 V_hig
+ 7.910010000e-07 V_hig
+ 7.911000000e-07 V_hig
+ 7.911010000e-07 V_hig
+ 7.912000000e-07 V_hig
+ 7.912010000e-07 V_hig
+ 7.913000000e-07 V_hig
+ 7.913010000e-07 V_hig
+ 7.914000000e-07 V_hig
+ 7.914010000e-07 V_hig
+ 7.915000000e-07 V_hig
+ 7.915010000e-07 V_hig
+ 7.916000000e-07 V_hig
+ 7.916010000e-07 V_hig
+ 7.917000000e-07 V_hig
+ 7.917010000e-07 V_hig
+ 7.918000000e-07 V_hig
+ 7.918010000e-07 V_hig
+ 7.919000000e-07 V_hig
+ 7.919010000e-07 V_low
+ 7.920000000e-07 V_low
+ 7.920010000e-07 V_low
+ 7.921000000e-07 V_low
+ 7.921010000e-07 V_low
+ 7.922000000e-07 V_low
+ 7.922010000e-07 V_low
+ 7.923000000e-07 V_low
+ 7.923010000e-07 V_low
+ 7.924000000e-07 V_low
+ 7.924010000e-07 V_low
+ 7.925000000e-07 V_low
+ 7.925010000e-07 V_low
+ 7.926000000e-07 V_low
+ 7.926010000e-07 V_low
+ 7.927000000e-07 V_low
+ 7.927010000e-07 V_low
+ 7.928000000e-07 V_low
+ 7.928010000e-07 V_low
+ 7.929000000e-07 V_low
+ 7.929010000e-07 V_hig
+ 7.930000000e-07 V_hig
+ 7.930010000e-07 V_hig
+ 7.931000000e-07 V_hig
+ 7.931010000e-07 V_hig
+ 7.932000000e-07 V_hig
+ 7.932010000e-07 V_hig
+ 7.933000000e-07 V_hig
+ 7.933010000e-07 V_hig
+ 7.934000000e-07 V_hig
+ 7.934010000e-07 V_hig
+ 7.935000000e-07 V_hig
+ 7.935010000e-07 V_hig
+ 7.936000000e-07 V_hig
+ 7.936010000e-07 V_hig
+ 7.937000000e-07 V_hig
+ 7.937010000e-07 V_hig
+ 7.938000000e-07 V_hig
+ 7.938010000e-07 V_hig
+ 7.939000000e-07 V_hig
+ 7.939010000e-07 V_low
+ 7.940000000e-07 V_low
+ 7.940010000e-07 V_low
+ 7.941000000e-07 V_low
+ 7.941010000e-07 V_low
+ 7.942000000e-07 V_low
+ 7.942010000e-07 V_low
+ 7.943000000e-07 V_low
+ 7.943010000e-07 V_low
+ 7.944000000e-07 V_low
+ 7.944010000e-07 V_low
+ 7.945000000e-07 V_low
+ 7.945010000e-07 V_low
+ 7.946000000e-07 V_low
+ 7.946010000e-07 V_low
+ 7.947000000e-07 V_low
+ 7.947010000e-07 V_low
+ 7.948000000e-07 V_low
+ 7.948010000e-07 V_low
+ 7.949000000e-07 V_low
+ 7.949010000e-07 V_hig
+ 7.950000000e-07 V_hig
+ 7.950010000e-07 V_hig
+ 7.951000000e-07 V_hig
+ 7.951010000e-07 V_hig
+ 7.952000000e-07 V_hig
+ 7.952010000e-07 V_hig
+ 7.953000000e-07 V_hig
+ 7.953010000e-07 V_hig
+ 7.954000000e-07 V_hig
+ 7.954010000e-07 V_hig
+ 7.955000000e-07 V_hig
+ 7.955010000e-07 V_hig
+ 7.956000000e-07 V_hig
+ 7.956010000e-07 V_hig
+ 7.957000000e-07 V_hig
+ 7.957010000e-07 V_hig
+ 7.958000000e-07 V_hig
+ 7.958010000e-07 V_hig
+ 7.959000000e-07 V_hig
+ 7.959010000e-07 V_low
+ 7.960000000e-07 V_low
+ 7.960010000e-07 V_low
+ 7.961000000e-07 V_low
+ 7.961010000e-07 V_low
+ 7.962000000e-07 V_low
+ 7.962010000e-07 V_low
+ 7.963000000e-07 V_low
+ 7.963010000e-07 V_low
+ 7.964000000e-07 V_low
+ 7.964010000e-07 V_low
+ 7.965000000e-07 V_low
+ 7.965010000e-07 V_low
+ 7.966000000e-07 V_low
+ 7.966010000e-07 V_low
+ 7.967000000e-07 V_low
+ 7.967010000e-07 V_low
+ 7.968000000e-07 V_low
+ 7.968010000e-07 V_low
+ 7.969000000e-07 V_low
+ 7.969010000e-07 V_low
+ 7.970000000e-07 V_low
+ 7.970010000e-07 V_low
+ 7.971000000e-07 V_low
+ 7.971010000e-07 V_low
+ 7.972000000e-07 V_low
+ 7.972010000e-07 V_low
+ 7.973000000e-07 V_low
+ 7.973010000e-07 V_low
+ 7.974000000e-07 V_low
+ 7.974010000e-07 V_low
+ 7.975000000e-07 V_low
+ 7.975010000e-07 V_low
+ 7.976000000e-07 V_low
+ 7.976010000e-07 V_low
+ 7.977000000e-07 V_low
+ 7.977010000e-07 V_low
+ 7.978000000e-07 V_low
+ 7.978010000e-07 V_low
+ 7.979000000e-07 V_low
+ 7.979010000e-07 V_hig
+ 7.980000000e-07 V_hig
+ 7.980010000e-07 V_hig
+ 7.981000000e-07 V_hig
+ 7.981010000e-07 V_hig
+ 7.982000000e-07 V_hig
+ 7.982010000e-07 V_hig
+ 7.983000000e-07 V_hig
+ 7.983010000e-07 V_hig
+ 7.984000000e-07 V_hig
+ 7.984010000e-07 V_hig
+ 7.985000000e-07 V_hig
+ 7.985010000e-07 V_hig
+ 7.986000000e-07 V_hig
+ 7.986010000e-07 V_hig
+ 7.987000000e-07 V_hig
+ 7.987010000e-07 V_hig
+ 7.988000000e-07 V_hig
+ 7.988010000e-07 V_hig
+ 7.989000000e-07 V_hig
+ 7.989010000e-07 V_low
+ 7.990000000e-07 V_low
+ 7.990010000e-07 V_low
+ 7.991000000e-07 V_low
+ 7.991010000e-07 V_low
+ 7.992000000e-07 V_low
+ 7.992010000e-07 V_low
+ 7.993000000e-07 V_low
+ 7.993010000e-07 V_low
+ 7.994000000e-07 V_low
+ 7.994010000e-07 V_low
+ 7.995000000e-07 V_low
+ 7.995010000e-07 V_low
+ 7.996000000e-07 V_low
+ 7.996010000e-07 V_low
+ 7.997000000e-07 V_low
+ 7.997010000e-07 V_low
+ 7.998000000e-07 V_low
+ 7.998010000e-07 V_low
+ 7.999000000e-07 V_low
+ 7.999010000e-07 V_hig
+ 8.000000000e-07 V_hig
+ 8.000010000e-07 V_hig
+ 8.001000000e-07 V_hig
+ 8.001010000e-07 V_hig
+ 8.002000000e-07 V_hig
+ 8.002010000e-07 V_hig
+ 8.003000000e-07 V_hig
+ 8.003010000e-07 V_hig
+ 8.004000000e-07 V_hig
+ 8.004010000e-07 V_hig
+ 8.005000000e-07 V_hig
+ 8.005010000e-07 V_hig
+ 8.006000000e-07 V_hig
+ 8.006010000e-07 V_hig
+ 8.007000000e-07 V_hig
+ 8.007010000e-07 V_hig
+ 8.008000000e-07 V_hig
+ 8.008010000e-07 V_hig
+ 8.009000000e-07 V_hig
+ 8.009010000e-07 V_hig
+ 8.010000000e-07 V_hig
+ 8.010010000e-07 V_hig
+ 8.011000000e-07 V_hig
+ 8.011010000e-07 V_hig
+ 8.012000000e-07 V_hig
+ 8.012010000e-07 V_hig
+ 8.013000000e-07 V_hig
+ 8.013010000e-07 V_hig
+ 8.014000000e-07 V_hig
+ 8.014010000e-07 V_hig
+ 8.015000000e-07 V_hig
+ 8.015010000e-07 V_hig
+ 8.016000000e-07 V_hig
+ 8.016010000e-07 V_hig
+ 8.017000000e-07 V_hig
+ 8.017010000e-07 V_hig
+ 8.018000000e-07 V_hig
+ 8.018010000e-07 V_hig
+ 8.019000000e-07 V_hig
+ 8.019010000e-07 V_low
+ 8.020000000e-07 V_low
+ 8.020010000e-07 V_low
+ 8.021000000e-07 V_low
+ 8.021010000e-07 V_low
+ 8.022000000e-07 V_low
+ 8.022010000e-07 V_low
+ 8.023000000e-07 V_low
+ 8.023010000e-07 V_low
+ 8.024000000e-07 V_low
+ 8.024010000e-07 V_low
+ 8.025000000e-07 V_low
+ 8.025010000e-07 V_low
+ 8.026000000e-07 V_low
+ 8.026010000e-07 V_low
+ 8.027000000e-07 V_low
+ 8.027010000e-07 V_low
+ 8.028000000e-07 V_low
+ 8.028010000e-07 V_low
+ 8.029000000e-07 V_low
+ 8.029010000e-07 V_hig
+ 8.030000000e-07 V_hig
+ 8.030010000e-07 V_hig
+ 8.031000000e-07 V_hig
+ 8.031010000e-07 V_hig
+ 8.032000000e-07 V_hig
+ 8.032010000e-07 V_hig
+ 8.033000000e-07 V_hig
+ 8.033010000e-07 V_hig
+ 8.034000000e-07 V_hig
+ 8.034010000e-07 V_hig
+ 8.035000000e-07 V_hig
+ 8.035010000e-07 V_hig
+ 8.036000000e-07 V_hig
+ 8.036010000e-07 V_hig
+ 8.037000000e-07 V_hig
+ 8.037010000e-07 V_hig
+ 8.038000000e-07 V_hig
+ 8.038010000e-07 V_hig
+ 8.039000000e-07 V_hig
+ 8.039010000e-07 V_low
+ 8.040000000e-07 V_low
+ 8.040010000e-07 V_low
+ 8.041000000e-07 V_low
+ 8.041010000e-07 V_low
+ 8.042000000e-07 V_low
+ 8.042010000e-07 V_low
+ 8.043000000e-07 V_low
+ 8.043010000e-07 V_low
+ 8.044000000e-07 V_low
+ 8.044010000e-07 V_low
+ 8.045000000e-07 V_low
+ 8.045010000e-07 V_low
+ 8.046000000e-07 V_low
+ 8.046010000e-07 V_low
+ 8.047000000e-07 V_low
+ 8.047010000e-07 V_low
+ 8.048000000e-07 V_low
+ 8.048010000e-07 V_low
+ 8.049000000e-07 V_low
+ 8.049010000e-07 V_hig
+ 8.050000000e-07 V_hig
+ 8.050010000e-07 V_hig
+ 8.051000000e-07 V_hig
+ 8.051010000e-07 V_hig
+ 8.052000000e-07 V_hig
+ 8.052010000e-07 V_hig
+ 8.053000000e-07 V_hig
+ 8.053010000e-07 V_hig
+ 8.054000000e-07 V_hig
+ 8.054010000e-07 V_hig
+ 8.055000000e-07 V_hig
+ 8.055010000e-07 V_hig
+ 8.056000000e-07 V_hig
+ 8.056010000e-07 V_hig
+ 8.057000000e-07 V_hig
+ 8.057010000e-07 V_hig
+ 8.058000000e-07 V_hig
+ 8.058010000e-07 V_hig
+ 8.059000000e-07 V_hig
+ 8.059010000e-07 V_low
+ 8.060000000e-07 V_low
+ 8.060010000e-07 V_low
+ 8.061000000e-07 V_low
+ 8.061010000e-07 V_low
+ 8.062000000e-07 V_low
+ 8.062010000e-07 V_low
+ 8.063000000e-07 V_low
+ 8.063010000e-07 V_low
+ 8.064000000e-07 V_low
+ 8.064010000e-07 V_low
+ 8.065000000e-07 V_low
+ 8.065010000e-07 V_low
+ 8.066000000e-07 V_low
+ 8.066010000e-07 V_low
+ 8.067000000e-07 V_low
+ 8.067010000e-07 V_low
+ 8.068000000e-07 V_low
+ 8.068010000e-07 V_low
+ 8.069000000e-07 V_low
+ 8.069010000e-07 V_hig
+ 8.070000000e-07 V_hig
+ 8.070010000e-07 V_hig
+ 8.071000000e-07 V_hig
+ 8.071010000e-07 V_hig
+ 8.072000000e-07 V_hig
+ 8.072010000e-07 V_hig
+ 8.073000000e-07 V_hig
+ 8.073010000e-07 V_hig
+ 8.074000000e-07 V_hig
+ 8.074010000e-07 V_hig
+ 8.075000000e-07 V_hig
+ 8.075010000e-07 V_hig
+ 8.076000000e-07 V_hig
+ 8.076010000e-07 V_hig
+ 8.077000000e-07 V_hig
+ 8.077010000e-07 V_hig
+ 8.078000000e-07 V_hig
+ 8.078010000e-07 V_hig
+ 8.079000000e-07 V_hig
+ 8.079010000e-07 V_low
+ 8.080000000e-07 V_low
+ 8.080010000e-07 V_low
+ 8.081000000e-07 V_low
+ 8.081010000e-07 V_low
+ 8.082000000e-07 V_low
+ 8.082010000e-07 V_low
+ 8.083000000e-07 V_low
+ 8.083010000e-07 V_low
+ 8.084000000e-07 V_low
+ 8.084010000e-07 V_low
+ 8.085000000e-07 V_low
+ 8.085010000e-07 V_low
+ 8.086000000e-07 V_low
+ 8.086010000e-07 V_low
+ 8.087000000e-07 V_low
+ 8.087010000e-07 V_low
+ 8.088000000e-07 V_low
+ 8.088010000e-07 V_low
+ 8.089000000e-07 V_low
+ 8.089010000e-07 V_low
+ 8.090000000e-07 V_low
+ 8.090010000e-07 V_low
+ 8.091000000e-07 V_low
+ 8.091010000e-07 V_low
+ 8.092000000e-07 V_low
+ 8.092010000e-07 V_low
+ 8.093000000e-07 V_low
+ 8.093010000e-07 V_low
+ 8.094000000e-07 V_low
+ 8.094010000e-07 V_low
+ 8.095000000e-07 V_low
+ 8.095010000e-07 V_low
+ 8.096000000e-07 V_low
+ 8.096010000e-07 V_low
+ 8.097000000e-07 V_low
+ 8.097010000e-07 V_low
+ 8.098000000e-07 V_low
+ 8.098010000e-07 V_low
+ 8.099000000e-07 V_low
+ 8.099010000e-07 V_hig
+ 8.100000000e-07 V_hig
+ 8.100010000e-07 V_hig
+ 8.101000000e-07 V_hig
+ 8.101010000e-07 V_hig
+ 8.102000000e-07 V_hig
+ 8.102010000e-07 V_hig
+ 8.103000000e-07 V_hig
+ 8.103010000e-07 V_hig
+ 8.104000000e-07 V_hig
+ 8.104010000e-07 V_hig
+ 8.105000000e-07 V_hig
+ 8.105010000e-07 V_hig
+ 8.106000000e-07 V_hig
+ 8.106010000e-07 V_hig
+ 8.107000000e-07 V_hig
+ 8.107010000e-07 V_hig
+ 8.108000000e-07 V_hig
+ 8.108010000e-07 V_hig
+ 8.109000000e-07 V_hig
+ 8.109010000e-07 V_low
+ 8.110000000e-07 V_low
+ 8.110010000e-07 V_low
+ 8.111000000e-07 V_low
+ 8.111010000e-07 V_low
+ 8.112000000e-07 V_low
+ 8.112010000e-07 V_low
+ 8.113000000e-07 V_low
+ 8.113010000e-07 V_low
+ 8.114000000e-07 V_low
+ 8.114010000e-07 V_low
+ 8.115000000e-07 V_low
+ 8.115010000e-07 V_low
+ 8.116000000e-07 V_low
+ 8.116010000e-07 V_low
+ 8.117000000e-07 V_low
+ 8.117010000e-07 V_low
+ 8.118000000e-07 V_low
+ 8.118010000e-07 V_low
+ 8.119000000e-07 V_low
+ 8.119010000e-07 V_low
+ 8.120000000e-07 V_low
+ 8.120010000e-07 V_low
+ 8.121000000e-07 V_low
+ 8.121010000e-07 V_low
+ 8.122000000e-07 V_low
+ 8.122010000e-07 V_low
+ 8.123000000e-07 V_low
+ 8.123010000e-07 V_low
+ 8.124000000e-07 V_low
+ 8.124010000e-07 V_low
+ 8.125000000e-07 V_low
+ 8.125010000e-07 V_low
+ 8.126000000e-07 V_low
+ 8.126010000e-07 V_low
+ 8.127000000e-07 V_low
+ 8.127010000e-07 V_low
+ 8.128000000e-07 V_low
+ 8.128010000e-07 V_low
+ 8.129000000e-07 V_low
+ 8.129010000e-07 V_low
+ 8.130000000e-07 V_low
+ 8.130010000e-07 V_low
+ 8.131000000e-07 V_low
+ 8.131010000e-07 V_low
+ 8.132000000e-07 V_low
+ 8.132010000e-07 V_low
+ 8.133000000e-07 V_low
+ 8.133010000e-07 V_low
+ 8.134000000e-07 V_low
+ 8.134010000e-07 V_low
+ 8.135000000e-07 V_low
+ 8.135010000e-07 V_low
+ 8.136000000e-07 V_low
+ 8.136010000e-07 V_low
+ 8.137000000e-07 V_low
+ 8.137010000e-07 V_low
+ 8.138000000e-07 V_low
+ 8.138010000e-07 V_low
+ 8.139000000e-07 V_low
+ 8.139010000e-07 V_hig
+ 8.140000000e-07 V_hig
+ 8.140010000e-07 V_hig
+ 8.141000000e-07 V_hig
+ 8.141010000e-07 V_hig
+ 8.142000000e-07 V_hig
+ 8.142010000e-07 V_hig
+ 8.143000000e-07 V_hig
+ 8.143010000e-07 V_hig
+ 8.144000000e-07 V_hig
+ 8.144010000e-07 V_hig
+ 8.145000000e-07 V_hig
+ 8.145010000e-07 V_hig
+ 8.146000000e-07 V_hig
+ 8.146010000e-07 V_hig
+ 8.147000000e-07 V_hig
+ 8.147010000e-07 V_hig
+ 8.148000000e-07 V_hig
+ 8.148010000e-07 V_hig
+ 8.149000000e-07 V_hig
+ 8.149010000e-07 V_hig
+ 8.150000000e-07 V_hig
+ 8.150010000e-07 V_hig
+ 8.151000000e-07 V_hig
+ 8.151010000e-07 V_hig
+ 8.152000000e-07 V_hig
+ 8.152010000e-07 V_hig
+ 8.153000000e-07 V_hig
+ 8.153010000e-07 V_hig
+ 8.154000000e-07 V_hig
+ 8.154010000e-07 V_hig
+ 8.155000000e-07 V_hig
+ 8.155010000e-07 V_hig
+ 8.156000000e-07 V_hig
+ 8.156010000e-07 V_hig
+ 8.157000000e-07 V_hig
+ 8.157010000e-07 V_hig
+ 8.158000000e-07 V_hig
+ 8.158010000e-07 V_hig
+ 8.159000000e-07 V_hig
+ 8.159010000e-07 V_hig
+ 8.160000000e-07 V_hig
+ 8.160010000e-07 V_hig
+ 8.161000000e-07 V_hig
+ 8.161010000e-07 V_hig
+ 8.162000000e-07 V_hig
+ 8.162010000e-07 V_hig
+ 8.163000000e-07 V_hig
+ 8.163010000e-07 V_hig
+ 8.164000000e-07 V_hig
+ 8.164010000e-07 V_hig
+ 8.165000000e-07 V_hig
+ 8.165010000e-07 V_hig
+ 8.166000000e-07 V_hig
+ 8.166010000e-07 V_hig
+ 8.167000000e-07 V_hig
+ 8.167010000e-07 V_hig
+ 8.168000000e-07 V_hig
+ 8.168010000e-07 V_hig
+ 8.169000000e-07 V_hig
+ 8.169010000e-07 V_hig
+ 8.170000000e-07 V_hig
+ 8.170010000e-07 V_hig
+ 8.171000000e-07 V_hig
+ 8.171010000e-07 V_hig
+ 8.172000000e-07 V_hig
+ 8.172010000e-07 V_hig
+ 8.173000000e-07 V_hig
+ 8.173010000e-07 V_hig
+ 8.174000000e-07 V_hig
+ 8.174010000e-07 V_hig
+ 8.175000000e-07 V_hig
+ 8.175010000e-07 V_hig
+ 8.176000000e-07 V_hig
+ 8.176010000e-07 V_hig
+ 8.177000000e-07 V_hig
+ 8.177010000e-07 V_hig
+ 8.178000000e-07 V_hig
+ 8.178010000e-07 V_hig
+ 8.179000000e-07 V_hig
+ 8.179010000e-07 V_hig
+ 8.180000000e-07 V_hig
+ 8.180010000e-07 V_hig
+ 8.181000000e-07 V_hig
+ 8.181010000e-07 V_hig
+ 8.182000000e-07 V_hig
+ 8.182010000e-07 V_hig
+ 8.183000000e-07 V_hig
+ 8.183010000e-07 V_hig
+ 8.184000000e-07 V_hig
+ 8.184010000e-07 V_hig
+ 8.185000000e-07 V_hig
+ 8.185010000e-07 V_hig
+ 8.186000000e-07 V_hig
+ 8.186010000e-07 V_hig
+ 8.187000000e-07 V_hig
+ 8.187010000e-07 V_hig
+ 8.188000000e-07 V_hig
+ 8.188010000e-07 V_hig
+ 8.189000000e-07 V_hig
+ 8.189010000e-07 V_low
+ 8.190000000e-07 V_low
+ 8.190010000e-07 V_low
+ 8.191000000e-07 V_low
+ 8.191010000e-07 V_low
+ 8.192000000e-07 V_low
+ 8.192010000e-07 V_low
+ 8.193000000e-07 V_low
+ 8.193010000e-07 V_low
+ 8.194000000e-07 V_low
+ 8.194010000e-07 V_low
+ 8.195000000e-07 V_low
+ 8.195010000e-07 V_low
+ 8.196000000e-07 V_low
+ 8.196010000e-07 V_low
+ 8.197000000e-07 V_low
+ 8.197010000e-07 V_low
+ 8.198000000e-07 V_low
+ 8.198010000e-07 V_low
+ 8.199000000e-07 V_low
+ 8.199010000e-07 V_hig
+ 8.200000000e-07 V_hig
+ 8.200010000e-07 V_hig
+ 8.201000000e-07 V_hig
+ 8.201010000e-07 V_hig
+ 8.202000000e-07 V_hig
+ 8.202010000e-07 V_hig
+ 8.203000000e-07 V_hig
+ 8.203010000e-07 V_hig
+ 8.204000000e-07 V_hig
+ 8.204010000e-07 V_hig
+ 8.205000000e-07 V_hig
+ 8.205010000e-07 V_hig
+ 8.206000000e-07 V_hig
+ 8.206010000e-07 V_hig
+ 8.207000000e-07 V_hig
+ 8.207010000e-07 V_hig
+ 8.208000000e-07 V_hig
+ 8.208010000e-07 V_hig
+ 8.209000000e-07 V_hig
+ 8.209010000e-07 V_hig
+ 8.210000000e-07 V_hig
+ 8.210010000e-07 V_hig
+ 8.211000000e-07 V_hig
+ 8.211010000e-07 V_hig
+ 8.212000000e-07 V_hig
+ 8.212010000e-07 V_hig
+ 8.213000000e-07 V_hig
+ 8.213010000e-07 V_hig
+ 8.214000000e-07 V_hig
+ 8.214010000e-07 V_hig
+ 8.215000000e-07 V_hig
+ 8.215010000e-07 V_hig
+ 8.216000000e-07 V_hig
+ 8.216010000e-07 V_hig
+ 8.217000000e-07 V_hig
+ 8.217010000e-07 V_hig
+ 8.218000000e-07 V_hig
+ 8.218010000e-07 V_hig
+ 8.219000000e-07 V_hig
+ 8.219010000e-07 V_hig
+ 8.220000000e-07 V_hig
+ 8.220010000e-07 V_hig
+ 8.221000000e-07 V_hig
+ 8.221010000e-07 V_hig
+ 8.222000000e-07 V_hig
+ 8.222010000e-07 V_hig
+ 8.223000000e-07 V_hig
+ 8.223010000e-07 V_hig
+ 8.224000000e-07 V_hig
+ 8.224010000e-07 V_hig
+ 8.225000000e-07 V_hig
+ 8.225010000e-07 V_hig
+ 8.226000000e-07 V_hig
+ 8.226010000e-07 V_hig
+ 8.227000000e-07 V_hig
+ 8.227010000e-07 V_hig
+ 8.228000000e-07 V_hig
+ 8.228010000e-07 V_hig
+ 8.229000000e-07 V_hig
+ 8.229010000e-07 V_hig
+ 8.230000000e-07 V_hig
+ 8.230010000e-07 V_hig
+ 8.231000000e-07 V_hig
+ 8.231010000e-07 V_hig
+ 8.232000000e-07 V_hig
+ 8.232010000e-07 V_hig
+ 8.233000000e-07 V_hig
+ 8.233010000e-07 V_hig
+ 8.234000000e-07 V_hig
+ 8.234010000e-07 V_hig
+ 8.235000000e-07 V_hig
+ 8.235010000e-07 V_hig
+ 8.236000000e-07 V_hig
+ 8.236010000e-07 V_hig
+ 8.237000000e-07 V_hig
+ 8.237010000e-07 V_hig
+ 8.238000000e-07 V_hig
+ 8.238010000e-07 V_hig
+ 8.239000000e-07 V_hig
+ 8.239010000e-07 V_hig
+ 8.240000000e-07 V_hig
+ 8.240010000e-07 V_hig
+ 8.241000000e-07 V_hig
+ 8.241010000e-07 V_hig
+ 8.242000000e-07 V_hig
+ 8.242010000e-07 V_hig
+ 8.243000000e-07 V_hig
+ 8.243010000e-07 V_hig
+ 8.244000000e-07 V_hig
+ 8.244010000e-07 V_hig
+ 8.245000000e-07 V_hig
+ 8.245010000e-07 V_hig
+ 8.246000000e-07 V_hig
+ 8.246010000e-07 V_hig
+ 8.247000000e-07 V_hig
+ 8.247010000e-07 V_hig
+ 8.248000000e-07 V_hig
+ 8.248010000e-07 V_hig
+ 8.249000000e-07 V_hig
+ 8.249010000e-07 V_low
+ 8.250000000e-07 V_low
+ 8.250010000e-07 V_low
+ 8.251000000e-07 V_low
+ 8.251010000e-07 V_low
+ 8.252000000e-07 V_low
+ 8.252010000e-07 V_low
+ 8.253000000e-07 V_low
+ 8.253010000e-07 V_low
+ 8.254000000e-07 V_low
+ 8.254010000e-07 V_low
+ 8.255000000e-07 V_low
+ 8.255010000e-07 V_low
+ 8.256000000e-07 V_low
+ 8.256010000e-07 V_low
+ 8.257000000e-07 V_low
+ 8.257010000e-07 V_low
+ 8.258000000e-07 V_low
+ 8.258010000e-07 V_low
+ 8.259000000e-07 V_low
+ 8.259010000e-07 V_low
+ 8.260000000e-07 V_low
+ 8.260010000e-07 V_low
+ 8.261000000e-07 V_low
+ 8.261010000e-07 V_low
+ 8.262000000e-07 V_low
+ 8.262010000e-07 V_low
+ 8.263000000e-07 V_low
+ 8.263010000e-07 V_low
+ 8.264000000e-07 V_low
+ 8.264010000e-07 V_low
+ 8.265000000e-07 V_low
+ 8.265010000e-07 V_low
+ 8.266000000e-07 V_low
+ 8.266010000e-07 V_low
+ 8.267000000e-07 V_low
+ 8.267010000e-07 V_low
+ 8.268000000e-07 V_low
+ 8.268010000e-07 V_low
+ 8.269000000e-07 V_low
+ 8.269010000e-07 V_low
+ 8.270000000e-07 V_low
+ 8.270010000e-07 V_low
+ 8.271000000e-07 V_low
+ 8.271010000e-07 V_low
+ 8.272000000e-07 V_low
+ 8.272010000e-07 V_low
+ 8.273000000e-07 V_low
+ 8.273010000e-07 V_low
+ 8.274000000e-07 V_low
+ 8.274010000e-07 V_low
+ 8.275000000e-07 V_low
+ 8.275010000e-07 V_low
+ 8.276000000e-07 V_low
+ 8.276010000e-07 V_low
+ 8.277000000e-07 V_low
+ 8.277010000e-07 V_low
+ 8.278000000e-07 V_low
+ 8.278010000e-07 V_low
+ 8.279000000e-07 V_low
+ 8.279010000e-07 V_low
+ 8.280000000e-07 V_low
+ 8.280010000e-07 V_low
+ 8.281000000e-07 V_low
+ 8.281010000e-07 V_low
+ 8.282000000e-07 V_low
+ 8.282010000e-07 V_low
+ 8.283000000e-07 V_low
+ 8.283010000e-07 V_low
+ 8.284000000e-07 V_low
+ 8.284010000e-07 V_low
+ 8.285000000e-07 V_low
+ 8.285010000e-07 V_low
+ 8.286000000e-07 V_low
+ 8.286010000e-07 V_low
+ 8.287000000e-07 V_low
+ 8.287010000e-07 V_low
+ 8.288000000e-07 V_low
+ 8.288010000e-07 V_low
+ 8.289000000e-07 V_low
+ 8.289010000e-07 V_hig
+ 8.290000000e-07 V_hig
+ 8.290010000e-07 V_hig
+ 8.291000000e-07 V_hig
+ 8.291010000e-07 V_hig
+ 8.292000000e-07 V_hig
+ 8.292010000e-07 V_hig
+ 8.293000000e-07 V_hig
+ 8.293010000e-07 V_hig
+ 8.294000000e-07 V_hig
+ 8.294010000e-07 V_hig
+ 8.295000000e-07 V_hig
+ 8.295010000e-07 V_hig
+ 8.296000000e-07 V_hig
+ 8.296010000e-07 V_hig
+ 8.297000000e-07 V_hig
+ 8.297010000e-07 V_hig
+ 8.298000000e-07 V_hig
+ 8.298010000e-07 V_hig
+ 8.299000000e-07 V_hig
+ 8.299010000e-07 V_low
+ 8.300000000e-07 V_low
+ 8.300010000e-07 V_low
+ 8.301000000e-07 V_low
+ 8.301010000e-07 V_low
+ 8.302000000e-07 V_low
+ 8.302010000e-07 V_low
+ 8.303000000e-07 V_low
+ 8.303010000e-07 V_low
+ 8.304000000e-07 V_low
+ 8.304010000e-07 V_low
+ 8.305000000e-07 V_low
+ 8.305010000e-07 V_low
+ 8.306000000e-07 V_low
+ 8.306010000e-07 V_low
+ 8.307000000e-07 V_low
+ 8.307010000e-07 V_low
+ 8.308000000e-07 V_low
+ 8.308010000e-07 V_low
+ 8.309000000e-07 V_low
+ 8.309010000e-07 V_hig
+ 8.310000000e-07 V_hig
+ 8.310010000e-07 V_hig
+ 8.311000000e-07 V_hig
+ 8.311010000e-07 V_hig
+ 8.312000000e-07 V_hig
+ 8.312010000e-07 V_hig
+ 8.313000000e-07 V_hig
+ 8.313010000e-07 V_hig
+ 8.314000000e-07 V_hig
+ 8.314010000e-07 V_hig
+ 8.315000000e-07 V_hig
+ 8.315010000e-07 V_hig
+ 8.316000000e-07 V_hig
+ 8.316010000e-07 V_hig
+ 8.317000000e-07 V_hig
+ 8.317010000e-07 V_hig
+ 8.318000000e-07 V_hig
+ 8.318010000e-07 V_hig
+ 8.319000000e-07 V_hig
+ 8.319010000e-07 V_low
+ 8.320000000e-07 V_low
+ 8.320010000e-07 V_low
+ 8.321000000e-07 V_low
+ 8.321010000e-07 V_low
+ 8.322000000e-07 V_low
+ 8.322010000e-07 V_low
+ 8.323000000e-07 V_low
+ 8.323010000e-07 V_low
+ 8.324000000e-07 V_low
+ 8.324010000e-07 V_low
+ 8.325000000e-07 V_low
+ 8.325010000e-07 V_low
+ 8.326000000e-07 V_low
+ 8.326010000e-07 V_low
+ 8.327000000e-07 V_low
+ 8.327010000e-07 V_low
+ 8.328000000e-07 V_low
+ 8.328010000e-07 V_low
+ 8.329000000e-07 V_low
+ 8.329010000e-07 V_low
+ 8.330000000e-07 V_low
+ 8.330010000e-07 V_low
+ 8.331000000e-07 V_low
+ 8.331010000e-07 V_low
+ 8.332000000e-07 V_low
+ 8.332010000e-07 V_low
+ 8.333000000e-07 V_low
+ 8.333010000e-07 V_low
+ 8.334000000e-07 V_low
+ 8.334010000e-07 V_low
+ 8.335000000e-07 V_low
+ 8.335010000e-07 V_low
+ 8.336000000e-07 V_low
+ 8.336010000e-07 V_low
+ 8.337000000e-07 V_low
+ 8.337010000e-07 V_low
+ 8.338000000e-07 V_low
+ 8.338010000e-07 V_low
+ 8.339000000e-07 V_low
+ 8.339010000e-07 V_low
+ 8.340000000e-07 V_low
+ 8.340010000e-07 V_low
+ 8.341000000e-07 V_low
+ 8.341010000e-07 V_low
+ 8.342000000e-07 V_low
+ 8.342010000e-07 V_low
+ 8.343000000e-07 V_low
+ 8.343010000e-07 V_low
+ 8.344000000e-07 V_low
+ 8.344010000e-07 V_low
+ 8.345000000e-07 V_low
+ 8.345010000e-07 V_low
+ 8.346000000e-07 V_low
+ 8.346010000e-07 V_low
+ 8.347000000e-07 V_low
+ 8.347010000e-07 V_low
+ 8.348000000e-07 V_low
+ 8.348010000e-07 V_low
+ 8.349000000e-07 V_low
+ 8.349010000e-07 V_low
+ 8.350000000e-07 V_low
+ 8.350010000e-07 V_low
+ 8.351000000e-07 V_low
+ 8.351010000e-07 V_low
+ 8.352000000e-07 V_low
+ 8.352010000e-07 V_low
+ 8.353000000e-07 V_low
+ 8.353010000e-07 V_low
+ 8.354000000e-07 V_low
+ 8.354010000e-07 V_low
+ 8.355000000e-07 V_low
+ 8.355010000e-07 V_low
+ 8.356000000e-07 V_low
+ 8.356010000e-07 V_low
+ 8.357000000e-07 V_low
+ 8.357010000e-07 V_low
+ 8.358000000e-07 V_low
+ 8.358010000e-07 V_low
+ 8.359000000e-07 V_low
+ 8.359010000e-07 V_hig
+ 8.360000000e-07 V_hig
+ 8.360010000e-07 V_hig
+ 8.361000000e-07 V_hig
+ 8.361010000e-07 V_hig
+ 8.362000000e-07 V_hig
+ 8.362010000e-07 V_hig
+ 8.363000000e-07 V_hig
+ 8.363010000e-07 V_hig
+ 8.364000000e-07 V_hig
+ 8.364010000e-07 V_hig
+ 8.365000000e-07 V_hig
+ 8.365010000e-07 V_hig
+ 8.366000000e-07 V_hig
+ 8.366010000e-07 V_hig
+ 8.367000000e-07 V_hig
+ 8.367010000e-07 V_hig
+ 8.368000000e-07 V_hig
+ 8.368010000e-07 V_hig
+ 8.369000000e-07 V_hig
+ 8.369010000e-07 V_low
+ 8.370000000e-07 V_low
+ 8.370010000e-07 V_low
+ 8.371000000e-07 V_low
+ 8.371010000e-07 V_low
+ 8.372000000e-07 V_low
+ 8.372010000e-07 V_low
+ 8.373000000e-07 V_low
+ 8.373010000e-07 V_low
+ 8.374000000e-07 V_low
+ 8.374010000e-07 V_low
+ 8.375000000e-07 V_low
+ 8.375010000e-07 V_low
+ 8.376000000e-07 V_low
+ 8.376010000e-07 V_low
+ 8.377000000e-07 V_low
+ 8.377010000e-07 V_low
+ 8.378000000e-07 V_low
+ 8.378010000e-07 V_low
+ 8.379000000e-07 V_low
+ 8.379010000e-07 V_low
+ 8.380000000e-07 V_low
+ 8.380010000e-07 V_low
+ 8.381000000e-07 V_low
+ 8.381010000e-07 V_low
+ 8.382000000e-07 V_low
+ 8.382010000e-07 V_low
+ 8.383000000e-07 V_low
+ 8.383010000e-07 V_low
+ 8.384000000e-07 V_low
+ 8.384010000e-07 V_low
+ 8.385000000e-07 V_low
+ 8.385010000e-07 V_low
+ 8.386000000e-07 V_low
+ 8.386010000e-07 V_low
+ 8.387000000e-07 V_low
+ 8.387010000e-07 V_low
+ 8.388000000e-07 V_low
+ 8.388010000e-07 V_low
+ 8.389000000e-07 V_low
+ 8.389010000e-07 V_hig
+ 8.390000000e-07 V_hig
+ 8.390010000e-07 V_hig
+ 8.391000000e-07 V_hig
+ 8.391010000e-07 V_hig
+ 8.392000000e-07 V_hig
+ 8.392010000e-07 V_hig
+ 8.393000000e-07 V_hig
+ 8.393010000e-07 V_hig
+ 8.394000000e-07 V_hig
+ 8.394010000e-07 V_hig
+ 8.395000000e-07 V_hig
+ 8.395010000e-07 V_hig
+ 8.396000000e-07 V_hig
+ 8.396010000e-07 V_hig
+ 8.397000000e-07 V_hig
+ 8.397010000e-07 V_hig
+ 8.398000000e-07 V_hig
+ 8.398010000e-07 V_hig
+ 8.399000000e-07 V_hig
+ 8.399010000e-07 V_hig
+ 8.400000000e-07 V_hig
+ 8.400010000e-07 V_hig
+ 8.401000000e-07 V_hig
+ 8.401010000e-07 V_hig
+ 8.402000000e-07 V_hig
+ 8.402010000e-07 V_hig
+ 8.403000000e-07 V_hig
+ 8.403010000e-07 V_hig
+ 8.404000000e-07 V_hig
+ 8.404010000e-07 V_hig
+ 8.405000000e-07 V_hig
+ 8.405010000e-07 V_hig
+ 8.406000000e-07 V_hig
+ 8.406010000e-07 V_hig
+ 8.407000000e-07 V_hig
+ 8.407010000e-07 V_hig
+ 8.408000000e-07 V_hig
+ 8.408010000e-07 V_hig
+ 8.409000000e-07 V_hig
+ 8.409010000e-07 V_low
+ 8.410000000e-07 V_low
+ 8.410010000e-07 V_low
+ 8.411000000e-07 V_low
+ 8.411010000e-07 V_low
+ 8.412000000e-07 V_low
+ 8.412010000e-07 V_low
+ 8.413000000e-07 V_low
+ 8.413010000e-07 V_low
+ 8.414000000e-07 V_low
+ 8.414010000e-07 V_low
+ 8.415000000e-07 V_low
+ 8.415010000e-07 V_low
+ 8.416000000e-07 V_low
+ 8.416010000e-07 V_low
+ 8.417000000e-07 V_low
+ 8.417010000e-07 V_low
+ 8.418000000e-07 V_low
+ 8.418010000e-07 V_low
+ 8.419000000e-07 V_low
+ 8.419010000e-07 V_low
+ 8.420000000e-07 V_low
+ 8.420010000e-07 V_low
+ 8.421000000e-07 V_low
+ 8.421010000e-07 V_low
+ 8.422000000e-07 V_low
+ 8.422010000e-07 V_low
+ 8.423000000e-07 V_low
+ 8.423010000e-07 V_low
+ 8.424000000e-07 V_low
+ 8.424010000e-07 V_low
+ 8.425000000e-07 V_low
+ 8.425010000e-07 V_low
+ 8.426000000e-07 V_low
+ 8.426010000e-07 V_low
+ 8.427000000e-07 V_low
+ 8.427010000e-07 V_low
+ 8.428000000e-07 V_low
+ 8.428010000e-07 V_low
+ 8.429000000e-07 V_low
+ 8.429010000e-07 V_hig
+ 8.430000000e-07 V_hig
+ 8.430010000e-07 V_hig
+ 8.431000000e-07 V_hig
+ 8.431010000e-07 V_hig
+ 8.432000000e-07 V_hig
+ 8.432010000e-07 V_hig
+ 8.433000000e-07 V_hig
+ 8.433010000e-07 V_hig
+ 8.434000000e-07 V_hig
+ 8.434010000e-07 V_hig
+ 8.435000000e-07 V_hig
+ 8.435010000e-07 V_hig
+ 8.436000000e-07 V_hig
+ 8.436010000e-07 V_hig
+ 8.437000000e-07 V_hig
+ 8.437010000e-07 V_hig
+ 8.438000000e-07 V_hig
+ 8.438010000e-07 V_hig
+ 8.439000000e-07 V_hig
+ 8.439010000e-07 V_hig
+ 8.440000000e-07 V_hig
+ 8.440010000e-07 V_hig
+ 8.441000000e-07 V_hig
+ 8.441010000e-07 V_hig
+ 8.442000000e-07 V_hig
+ 8.442010000e-07 V_hig
+ 8.443000000e-07 V_hig
+ 8.443010000e-07 V_hig
+ 8.444000000e-07 V_hig
+ 8.444010000e-07 V_hig
+ 8.445000000e-07 V_hig
+ 8.445010000e-07 V_hig
+ 8.446000000e-07 V_hig
+ 8.446010000e-07 V_hig
+ 8.447000000e-07 V_hig
+ 8.447010000e-07 V_hig
+ 8.448000000e-07 V_hig
+ 8.448010000e-07 V_hig
+ 8.449000000e-07 V_hig
+ 8.449010000e-07 V_low
+ 8.450000000e-07 V_low
+ 8.450010000e-07 V_low
+ 8.451000000e-07 V_low
+ 8.451010000e-07 V_low
+ 8.452000000e-07 V_low
+ 8.452010000e-07 V_low
+ 8.453000000e-07 V_low
+ 8.453010000e-07 V_low
+ 8.454000000e-07 V_low
+ 8.454010000e-07 V_low
+ 8.455000000e-07 V_low
+ 8.455010000e-07 V_low
+ 8.456000000e-07 V_low
+ 8.456010000e-07 V_low
+ 8.457000000e-07 V_low
+ 8.457010000e-07 V_low
+ 8.458000000e-07 V_low
+ 8.458010000e-07 V_low
+ 8.459000000e-07 V_low
+ 8.459010000e-07 V_hig
+ 8.460000000e-07 V_hig
+ 8.460010000e-07 V_hig
+ 8.461000000e-07 V_hig
+ 8.461010000e-07 V_hig
+ 8.462000000e-07 V_hig
+ 8.462010000e-07 V_hig
+ 8.463000000e-07 V_hig
+ 8.463010000e-07 V_hig
+ 8.464000000e-07 V_hig
+ 8.464010000e-07 V_hig
+ 8.465000000e-07 V_hig
+ 8.465010000e-07 V_hig
+ 8.466000000e-07 V_hig
+ 8.466010000e-07 V_hig
+ 8.467000000e-07 V_hig
+ 8.467010000e-07 V_hig
+ 8.468000000e-07 V_hig
+ 8.468010000e-07 V_hig
+ 8.469000000e-07 V_hig
+ 8.469010000e-07 V_hig
+ 8.470000000e-07 V_hig
+ 8.470010000e-07 V_hig
+ 8.471000000e-07 V_hig
+ 8.471010000e-07 V_hig
+ 8.472000000e-07 V_hig
+ 8.472010000e-07 V_hig
+ 8.473000000e-07 V_hig
+ 8.473010000e-07 V_hig
+ 8.474000000e-07 V_hig
+ 8.474010000e-07 V_hig
+ 8.475000000e-07 V_hig
+ 8.475010000e-07 V_hig
+ 8.476000000e-07 V_hig
+ 8.476010000e-07 V_hig
+ 8.477000000e-07 V_hig
+ 8.477010000e-07 V_hig
+ 8.478000000e-07 V_hig
+ 8.478010000e-07 V_hig
+ 8.479000000e-07 V_hig
+ 8.479010000e-07 V_hig
+ 8.480000000e-07 V_hig
+ 8.480010000e-07 V_hig
+ 8.481000000e-07 V_hig
+ 8.481010000e-07 V_hig
+ 8.482000000e-07 V_hig
+ 8.482010000e-07 V_hig
+ 8.483000000e-07 V_hig
+ 8.483010000e-07 V_hig
+ 8.484000000e-07 V_hig
+ 8.484010000e-07 V_hig
+ 8.485000000e-07 V_hig
+ 8.485010000e-07 V_hig
+ 8.486000000e-07 V_hig
+ 8.486010000e-07 V_hig
+ 8.487000000e-07 V_hig
+ 8.487010000e-07 V_hig
+ 8.488000000e-07 V_hig
+ 8.488010000e-07 V_hig
+ 8.489000000e-07 V_hig
+ 8.489010000e-07 V_low
+ 8.490000000e-07 V_low
+ 8.490010000e-07 V_low
+ 8.491000000e-07 V_low
+ 8.491010000e-07 V_low
+ 8.492000000e-07 V_low
+ 8.492010000e-07 V_low
+ 8.493000000e-07 V_low
+ 8.493010000e-07 V_low
+ 8.494000000e-07 V_low
+ 8.494010000e-07 V_low
+ 8.495000000e-07 V_low
+ 8.495010000e-07 V_low
+ 8.496000000e-07 V_low
+ 8.496010000e-07 V_low
+ 8.497000000e-07 V_low
+ 8.497010000e-07 V_low
+ 8.498000000e-07 V_low
+ 8.498010000e-07 V_low
+ 8.499000000e-07 V_low
+ 8.499010000e-07 V_low
+ 8.500000000e-07 V_low
+ 8.500010000e-07 V_low
+ 8.501000000e-07 V_low
+ 8.501010000e-07 V_low
+ 8.502000000e-07 V_low
+ 8.502010000e-07 V_low
+ 8.503000000e-07 V_low
+ 8.503010000e-07 V_low
+ 8.504000000e-07 V_low
+ 8.504010000e-07 V_low
+ 8.505000000e-07 V_low
+ 8.505010000e-07 V_low
+ 8.506000000e-07 V_low
+ 8.506010000e-07 V_low
+ 8.507000000e-07 V_low
+ 8.507010000e-07 V_low
+ 8.508000000e-07 V_low
+ 8.508010000e-07 V_low
+ 8.509000000e-07 V_low
+ 8.509010000e-07 V_hig
+ 8.510000000e-07 V_hig
+ 8.510010000e-07 V_hig
+ 8.511000000e-07 V_hig
+ 8.511010000e-07 V_hig
+ 8.512000000e-07 V_hig
+ 8.512010000e-07 V_hig
+ 8.513000000e-07 V_hig
+ 8.513010000e-07 V_hig
+ 8.514000000e-07 V_hig
+ 8.514010000e-07 V_hig
+ 8.515000000e-07 V_hig
+ 8.515010000e-07 V_hig
+ 8.516000000e-07 V_hig
+ 8.516010000e-07 V_hig
+ 8.517000000e-07 V_hig
+ 8.517010000e-07 V_hig
+ 8.518000000e-07 V_hig
+ 8.518010000e-07 V_hig
+ 8.519000000e-07 V_hig
+ 8.519010000e-07 V_hig
+ 8.520000000e-07 V_hig
+ 8.520010000e-07 V_hig
+ 8.521000000e-07 V_hig
+ 8.521010000e-07 V_hig
+ 8.522000000e-07 V_hig
+ 8.522010000e-07 V_hig
+ 8.523000000e-07 V_hig
+ 8.523010000e-07 V_hig
+ 8.524000000e-07 V_hig
+ 8.524010000e-07 V_hig
+ 8.525000000e-07 V_hig
+ 8.525010000e-07 V_hig
+ 8.526000000e-07 V_hig
+ 8.526010000e-07 V_hig
+ 8.527000000e-07 V_hig
+ 8.527010000e-07 V_hig
+ 8.528000000e-07 V_hig
+ 8.528010000e-07 V_hig
+ 8.529000000e-07 V_hig
+ 8.529010000e-07 V_low
+ 8.530000000e-07 V_low
+ 8.530010000e-07 V_low
+ 8.531000000e-07 V_low
+ 8.531010000e-07 V_low
+ 8.532000000e-07 V_low
+ 8.532010000e-07 V_low
+ 8.533000000e-07 V_low
+ 8.533010000e-07 V_low
+ 8.534000000e-07 V_low
+ 8.534010000e-07 V_low
+ 8.535000000e-07 V_low
+ 8.535010000e-07 V_low
+ 8.536000000e-07 V_low
+ 8.536010000e-07 V_low
+ 8.537000000e-07 V_low
+ 8.537010000e-07 V_low
+ 8.538000000e-07 V_low
+ 8.538010000e-07 V_low
+ 8.539000000e-07 V_low
+ 8.539010000e-07 V_hig
+ 8.540000000e-07 V_hig
+ 8.540010000e-07 V_hig
+ 8.541000000e-07 V_hig
+ 8.541010000e-07 V_hig
+ 8.542000000e-07 V_hig
+ 8.542010000e-07 V_hig
+ 8.543000000e-07 V_hig
+ 8.543010000e-07 V_hig
+ 8.544000000e-07 V_hig
+ 8.544010000e-07 V_hig
+ 8.545000000e-07 V_hig
+ 8.545010000e-07 V_hig
+ 8.546000000e-07 V_hig
+ 8.546010000e-07 V_hig
+ 8.547000000e-07 V_hig
+ 8.547010000e-07 V_hig
+ 8.548000000e-07 V_hig
+ 8.548010000e-07 V_hig
+ 8.549000000e-07 V_hig
+ 8.549010000e-07 V_hig
+ 8.550000000e-07 V_hig
+ 8.550010000e-07 V_hig
+ 8.551000000e-07 V_hig
+ 8.551010000e-07 V_hig
+ 8.552000000e-07 V_hig
+ 8.552010000e-07 V_hig
+ 8.553000000e-07 V_hig
+ 8.553010000e-07 V_hig
+ 8.554000000e-07 V_hig
+ 8.554010000e-07 V_hig
+ 8.555000000e-07 V_hig
+ 8.555010000e-07 V_hig
+ 8.556000000e-07 V_hig
+ 8.556010000e-07 V_hig
+ 8.557000000e-07 V_hig
+ 8.557010000e-07 V_hig
+ 8.558000000e-07 V_hig
+ 8.558010000e-07 V_hig
+ 8.559000000e-07 V_hig
+ 8.559010000e-07 V_low
+ 8.560000000e-07 V_low
+ 8.560010000e-07 V_low
+ 8.561000000e-07 V_low
+ 8.561010000e-07 V_low
+ 8.562000000e-07 V_low
+ 8.562010000e-07 V_low
+ 8.563000000e-07 V_low
+ 8.563010000e-07 V_low
+ 8.564000000e-07 V_low
+ 8.564010000e-07 V_low
+ 8.565000000e-07 V_low
+ 8.565010000e-07 V_low
+ 8.566000000e-07 V_low
+ 8.566010000e-07 V_low
+ 8.567000000e-07 V_low
+ 8.567010000e-07 V_low
+ 8.568000000e-07 V_low
+ 8.568010000e-07 V_low
+ 8.569000000e-07 V_low
+ 8.569010000e-07 V_low
+ 8.570000000e-07 V_low
+ 8.570010000e-07 V_low
+ 8.571000000e-07 V_low
+ 8.571010000e-07 V_low
+ 8.572000000e-07 V_low
+ 8.572010000e-07 V_low
+ 8.573000000e-07 V_low
+ 8.573010000e-07 V_low
+ 8.574000000e-07 V_low
+ 8.574010000e-07 V_low
+ 8.575000000e-07 V_low
+ 8.575010000e-07 V_low
+ 8.576000000e-07 V_low
+ 8.576010000e-07 V_low
+ 8.577000000e-07 V_low
+ 8.577010000e-07 V_low
+ 8.578000000e-07 V_low
+ 8.578010000e-07 V_low
+ 8.579000000e-07 V_low
+ 8.579010000e-07 V_low
+ 8.580000000e-07 V_low
+ 8.580010000e-07 V_low
+ 8.581000000e-07 V_low
+ 8.581010000e-07 V_low
+ 8.582000000e-07 V_low
+ 8.582010000e-07 V_low
+ 8.583000000e-07 V_low
+ 8.583010000e-07 V_low
+ 8.584000000e-07 V_low
+ 8.584010000e-07 V_low
+ 8.585000000e-07 V_low
+ 8.585010000e-07 V_low
+ 8.586000000e-07 V_low
+ 8.586010000e-07 V_low
+ 8.587000000e-07 V_low
+ 8.587010000e-07 V_low
+ 8.588000000e-07 V_low
+ 8.588010000e-07 V_low
+ 8.589000000e-07 V_low
+ 8.589010000e-07 V_hig
+ 8.590000000e-07 V_hig
+ 8.590010000e-07 V_hig
+ 8.591000000e-07 V_hig
+ 8.591010000e-07 V_hig
+ 8.592000000e-07 V_hig
+ 8.592010000e-07 V_hig
+ 8.593000000e-07 V_hig
+ 8.593010000e-07 V_hig
+ 8.594000000e-07 V_hig
+ 8.594010000e-07 V_hig
+ 8.595000000e-07 V_hig
+ 8.595010000e-07 V_hig
+ 8.596000000e-07 V_hig
+ 8.596010000e-07 V_hig
+ 8.597000000e-07 V_hig
+ 8.597010000e-07 V_hig
+ 8.598000000e-07 V_hig
+ 8.598010000e-07 V_hig
+ 8.599000000e-07 V_hig
+ 8.599010000e-07 V_hig
+ 8.600000000e-07 V_hig
+ 8.600010000e-07 V_hig
+ 8.601000000e-07 V_hig
+ 8.601010000e-07 V_hig
+ 8.602000000e-07 V_hig
+ 8.602010000e-07 V_hig
+ 8.603000000e-07 V_hig
+ 8.603010000e-07 V_hig
+ 8.604000000e-07 V_hig
+ 8.604010000e-07 V_hig
+ 8.605000000e-07 V_hig
+ 8.605010000e-07 V_hig
+ 8.606000000e-07 V_hig
+ 8.606010000e-07 V_hig
+ 8.607000000e-07 V_hig
+ 8.607010000e-07 V_hig
+ 8.608000000e-07 V_hig
+ 8.608010000e-07 V_hig
+ 8.609000000e-07 V_hig
+ 8.609010000e-07 V_hig
+ 8.610000000e-07 V_hig
+ 8.610010000e-07 V_hig
+ 8.611000000e-07 V_hig
+ 8.611010000e-07 V_hig
+ 8.612000000e-07 V_hig
+ 8.612010000e-07 V_hig
+ 8.613000000e-07 V_hig
+ 8.613010000e-07 V_hig
+ 8.614000000e-07 V_hig
+ 8.614010000e-07 V_hig
+ 8.615000000e-07 V_hig
+ 8.615010000e-07 V_hig
+ 8.616000000e-07 V_hig
+ 8.616010000e-07 V_hig
+ 8.617000000e-07 V_hig
+ 8.617010000e-07 V_hig
+ 8.618000000e-07 V_hig
+ 8.618010000e-07 V_hig
+ 8.619000000e-07 V_hig
+ 8.619010000e-07 V_low
+ 8.620000000e-07 V_low
+ 8.620010000e-07 V_low
+ 8.621000000e-07 V_low
+ 8.621010000e-07 V_low
+ 8.622000000e-07 V_low
+ 8.622010000e-07 V_low
+ 8.623000000e-07 V_low
+ 8.623010000e-07 V_low
+ 8.624000000e-07 V_low
+ 8.624010000e-07 V_low
+ 8.625000000e-07 V_low
+ 8.625010000e-07 V_low
+ 8.626000000e-07 V_low
+ 8.626010000e-07 V_low
+ 8.627000000e-07 V_low
+ 8.627010000e-07 V_low
+ 8.628000000e-07 V_low
+ 8.628010000e-07 V_low
+ 8.629000000e-07 V_low
+ 8.629010000e-07 V_low
+ 8.630000000e-07 V_low
+ 8.630010000e-07 V_low
+ 8.631000000e-07 V_low
+ 8.631010000e-07 V_low
+ 8.632000000e-07 V_low
+ 8.632010000e-07 V_low
+ 8.633000000e-07 V_low
+ 8.633010000e-07 V_low
+ 8.634000000e-07 V_low
+ 8.634010000e-07 V_low
+ 8.635000000e-07 V_low
+ 8.635010000e-07 V_low
+ 8.636000000e-07 V_low
+ 8.636010000e-07 V_low
+ 8.637000000e-07 V_low
+ 8.637010000e-07 V_low
+ 8.638000000e-07 V_low
+ 8.638010000e-07 V_low
+ 8.639000000e-07 V_low
+ 8.639010000e-07 V_hig
+ 8.640000000e-07 V_hig
+ 8.640010000e-07 V_hig
+ 8.641000000e-07 V_hig
+ 8.641010000e-07 V_hig
+ 8.642000000e-07 V_hig
+ 8.642010000e-07 V_hig
+ 8.643000000e-07 V_hig
+ 8.643010000e-07 V_hig
+ 8.644000000e-07 V_hig
+ 8.644010000e-07 V_hig
+ 8.645000000e-07 V_hig
+ 8.645010000e-07 V_hig
+ 8.646000000e-07 V_hig
+ 8.646010000e-07 V_hig
+ 8.647000000e-07 V_hig
+ 8.647010000e-07 V_hig
+ 8.648000000e-07 V_hig
+ 8.648010000e-07 V_hig
+ 8.649000000e-07 V_hig
+ 8.649010000e-07 V_hig
+ 8.650000000e-07 V_hig
+ 8.650010000e-07 V_hig
+ 8.651000000e-07 V_hig
+ 8.651010000e-07 V_hig
+ 8.652000000e-07 V_hig
+ 8.652010000e-07 V_hig
+ 8.653000000e-07 V_hig
+ 8.653010000e-07 V_hig
+ 8.654000000e-07 V_hig
+ 8.654010000e-07 V_hig
+ 8.655000000e-07 V_hig
+ 8.655010000e-07 V_hig
+ 8.656000000e-07 V_hig
+ 8.656010000e-07 V_hig
+ 8.657000000e-07 V_hig
+ 8.657010000e-07 V_hig
+ 8.658000000e-07 V_hig
+ 8.658010000e-07 V_hig
+ 8.659000000e-07 V_hig
+ 8.659010000e-07 V_low
+ 8.660000000e-07 V_low
+ 8.660010000e-07 V_low
+ 8.661000000e-07 V_low
+ 8.661010000e-07 V_low
+ 8.662000000e-07 V_low
+ 8.662010000e-07 V_low
+ 8.663000000e-07 V_low
+ 8.663010000e-07 V_low
+ 8.664000000e-07 V_low
+ 8.664010000e-07 V_low
+ 8.665000000e-07 V_low
+ 8.665010000e-07 V_low
+ 8.666000000e-07 V_low
+ 8.666010000e-07 V_low
+ 8.667000000e-07 V_low
+ 8.667010000e-07 V_low
+ 8.668000000e-07 V_low
+ 8.668010000e-07 V_low
+ 8.669000000e-07 V_low
+ 8.669010000e-07 V_hig
+ 8.670000000e-07 V_hig
+ 8.670010000e-07 V_hig
+ 8.671000000e-07 V_hig
+ 8.671010000e-07 V_hig
+ 8.672000000e-07 V_hig
+ 8.672010000e-07 V_hig
+ 8.673000000e-07 V_hig
+ 8.673010000e-07 V_hig
+ 8.674000000e-07 V_hig
+ 8.674010000e-07 V_hig
+ 8.675000000e-07 V_hig
+ 8.675010000e-07 V_hig
+ 8.676000000e-07 V_hig
+ 8.676010000e-07 V_hig
+ 8.677000000e-07 V_hig
+ 8.677010000e-07 V_hig
+ 8.678000000e-07 V_hig
+ 8.678010000e-07 V_hig
+ 8.679000000e-07 V_hig
+ 8.679010000e-07 V_hig
+ 8.680000000e-07 V_hig
+ 8.680010000e-07 V_hig
+ 8.681000000e-07 V_hig
+ 8.681010000e-07 V_hig
+ 8.682000000e-07 V_hig
+ 8.682010000e-07 V_hig
+ 8.683000000e-07 V_hig
+ 8.683010000e-07 V_hig
+ 8.684000000e-07 V_hig
+ 8.684010000e-07 V_hig
+ 8.685000000e-07 V_hig
+ 8.685010000e-07 V_hig
+ 8.686000000e-07 V_hig
+ 8.686010000e-07 V_hig
+ 8.687000000e-07 V_hig
+ 8.687010000e-07 V_hig
+ 8.688000000e-07 V_hig
+ 8.688010000e-07 V_hig
+ 8.689000000e-07 V_hig
+ 8.689010000e-07 V_hig
+ 8.690000000e-07 V_hig
+ 8.690010000e-07 V_hig
+ 8.691000000e-07 V_hig
+ 8.691010000e-07 V_hig
+ 8.692000000e-07 V_hig
+ 8.692010000e-07 V_hig
+ 8.693000000e-07 V_hig
+ 8.693010000e-07 V_hig
+ 8.694000000e-07 V_hig
+ 8.694010000e-07 V_hig
+ 8.695000000e-07 V_hig
+ 8.695010000e-07 V_hig
+ 8.696000000e-07 V_hig
+ 8.696010000e-07 V_hig
+ 8.697000000e-07 V_hig
+ 8.697010000e-07 V_hig
+ 8.698000000e-07 V_hig
+ 8.698010000e-07 V_hig
+ 8.699000000e-07 V_hig
+ 8.699010000e-07 V_hig
+ 8.700000000e-07 V_hig
+ 8.700010000e-07 V_hig
+ 8.701000000e-07 V_hig
+ 8.701010000e-07 V_hig
+ 8.702000000e-07 V_hig
+ 8.702010000e-07 V_hig
+ 8.703000000e-07 V_hig
+ 8.703010000e-07 V_hig
+ 8.704000000e-07 V_hig
+ 8.704010000e-07 V_hig
+ 8.705000000e-07 V_hig
+ 8.705010000e-07 V_hig
+ 8.706000000e-07 V_hig
+ 8.706010000e-07 V_hig
+ 8.707000000e-07 V_hig
+ 8.707010000e-07 V_hig
+ 8.708000000e-07 V_hig
+ 8.708010000e-07 V_hig
+ 8.709000000e-07 V_hig
+ 8.709010000e-07 V_low
+ 8.710000000e-07 V_low
+ 8.710010000e-07 V_low
+ 8.711000000e-07 V_low
+ 8.711010000e-07 V_low
+ 8.712000000e-07 V_low
+ 8.712010000e-07 V_low
+ 8.713000000e-07 V_low
+ 8.713010000e-07 V_low
+ 8.714000000e-07 V_low
+ 8.714010000e-07 V_low
+ 8.715000000e-07 V_low
+ 8.715010000e-07 V_low
+ 8.716000000e-07 V_low
+ 8.716010000e-07 V_low
+ 8.717000000e-07 V_low
+ 8.717010000e-07 V_low
+ 8.718000000e-07 V_low
+ 8.718010000e-07 V_low
+ 8.719000000e-07 V_low
+ 8.719010000e-07 V_hig
+ 8.720000000e-07 V_hig
+ 8.720010000e-07 V_hig
+ 8.721000000e-07 V_hig
+ 8.721010000e-07 V_hig
+ 8.722000000e-07 V_hig
+ 8.722010000e-07 V_hig
+ 8.723000000e-07 V_hig
+ 8.723010000e-07 V_hig
+ 8.724000000e-07 V_hig
+ 8.724010000e-07 V_hig
+ 8.725000000e-07 V_hig
+ 8.725010000e-07 V_hig
+ 8.726000000e-07 V_hig
+ 8.726010000e-07 V_hig
+ 8.727000000e-07 V_hig
+ 8.727010000e-07 V_hig
+ 8.728000000e-07 V_hig
+ 8.728010000e-07 V_hig
+ 8.729000000e-07 V_hig
+ 8.729010000e-07 V_low
+ 8.730000000e-07 V_low
+ 8.730010000e-07 V_low
+ 8.731000000e-07 V_low
+ 8.731010000e-07 V_low
+ 8.732000000e-07 V_low
+ 8.732010000e-07 V_low
+ 8.733000000e-07 V_low
+ 8.733010000e-07 V_low
+ 8.734000000e-07 V_low
+ 8.734010000e-07 V_low
+ 8.735000000e-07 V_low
+ 8.735010000e-07 V_low
+ 8.736000000e-07 V_low
+ 8.736010000e-07 V_low
+ 8.737000000e-07 V_low
+ 8.737010000e-07 V_low
+ 8.738000000e-07 V_low
+ 8.738010000e-07 V_low
+ 8.739000000e-07 V_low
+ 8.739010000e-07 V_hig
+ 8.740000000e-07 V_hig
+ 8.740010000e-07 V_hig
+ 8.741000000e-07 V_hig
+ 8.741010000e-07 V_hig
+ 8.742000000e-07 V_hig
+ 8.742010000e-07 V_hig
+ 8.743000000e-07 V_hig
+ 8.743010000e-07 V_hig
+ 8.744000000e-07 V_hig
+ 8.744010000e-07 V_hig
+ 8.745000000e-07 V_hig
+ 8.745010000e-07 V_hig
+ 8.746000000e-07 V_hig
+ 8.746010000e-07 V_hig
+ 8.747000000e-07 V_hig
+ 8.747010000e-07 V_hig
+ 8.748000000e-07 V_hig
+ 8.748010000e-07 V_hig
+ 8.749000000e-07 V_hig
+ 8.749010000e-07 V_hig
+ 8.750000000e-07 V_hig
+ 8.750010000e-07 V_hig
+ 8.751000000e-07 V_hig
+ 8.751010000e-07 V_hig
+ 8.752000000e-07 V_hig
+ 8.752010000e-07 V_hig
+ 8.753000000e-07 V_hig
+ 8.753010000e-07 V_hig
+ 8.754000000e-07 V_hig
+ 8.754010000e-07 V_hig
+ 8.755000000e-07 V_hig
+ 8.755010000e-07 V_hig
+ 8.756000000e-07 V_hig
+ 8.756010000e-07 V_hig
+ 8.757000000e-07 V_hig
+ 8.757010000e-07 V_hig
+ 8.758000000e-07 V_hig
+ 8.758010000e-07 V_hig
+ 8.759000000e-07 V_hig
+ 8.759010000e-07 V_low
+ 8.760000000e-07 V_low
+ 8.760010000e-07 V_low
+ 8.761000000e-07 V_low
+ 8.761010000e-07 V_low
+ 8.762000000e-07 V_low
+ 8.762010000e-07 V_low
+ 8.763000000e-07 V_low
+ 8.763010000e-07 V_low
+ 8.764000000e-07 V_low
+ 8.764010000e-07 V_low
+ 8.765000000e-07 V_low
+ 8.765010000e-07 V_low
+ 8.766000000e-07 V_low
+ 8.766010000e-07 V_low
+ 8.767000000e-07 V_low
+ 8.767010000e-07 V_low
+ 8.768000000e-07 V_low
+ 8.768010000e-07 V_low
+ 8.769000000e-07 V_low
+ 8.769010000e-07 V_low
+ 8.770000000e-07 V_low
+ 8.770010000e-07 V_low
+ 8.771000000e-07 V_low
+ 8.771010000e-07 V_low
+ 8.772000000e-07 V_low
+ 8.772010000e-07 V_low
+ 8.773000000e-07 V_low
+ 8.773010000e-07 V_low
+ 8.774000000e-07 V_low
+ 8.774010000e-07 V_low
+ 8.775000000e-07 V_low
+ 8.775010000e-07 V_low
+ 8.776000000e-07 V_low
+ 8.776010000e-07 V_low
+ 8.777000000e-07 V_low
+ 8.777010000e-07 V_low
+ 8.778000000e-07 V_low
+ 8.778010000e-07 V_low
+ 8.779000000e-07 V_low
+ 8.779010000e-07 V_low
+ 8.780000000e-07 V_low
+ 8.780010000e-07 V_low
+ 8.781000000e-07 V_low
+ 8.781010000e-07 V_low
+ 8.782000000e-07 V_low
+ 8.782010000e-07 V_low
+ 8.783000000e-07 V_low
+ 8.783010000e-07 V_low
+ 8.784000000e-07 V_low
+ 8.784010000e-07 V_low
+ 8.785000000e-07 V_low
+ 8.785010000e-07 V_low
+ 8.786000000e-07 V_low
+ 8.786010000e-07 V_low
+ 8.787000000e-07 V_low
+ 8.787010000e-07 V_low
+ 8.788000000e-07 V_low
+ 8.788010000e-07 V_low
+ 8.789000000e-07 V_low
+ 8.789010000e-07 V_hig
+ 8.790000000e-07 V_hig
+ 8.790010000e-07 V_hig
+ 8.791000000e-07 V_hig
+ 8.791010000e-07 V_hig
+ 8.792000000e-07 V_hig
+ 8.792010000e-07 V_hig
+ 8.793000000e-07 V_hig
+ 8.793010000e-07 V_hig
+ 8.794000000e-07 V_hig
+ 8.794010000e-07 V_hig
+ 8.795000000e-07 V_hig
+ 8.795010000e-07 V_hig
+ 8.796000000e-07 V_hig
+ 8.796010000e-07 V_hig
+ 8.797000000e-07 V_hig
+ 8.797010000e-07 V_hig
+ 8.798000000e-07 V_hig
+ 8.798010000e-07 V_hig
+ 8.799000000e-07 V_hig
+ 8.799010000e-07 V_low
+ 8.800000000e-07 V_low
+ 8.800010000e-07 V_low
+ 8.801000000e-07 V_low
+ 8.801010000e-07 V_low
+ 8.802000000e-07 V_low
+ 8.802010000e-07 V_low
+ 8.803000000e-07 V_low
+ 8.803010000e-07 V_low
+ 8.804000000e-07 V_low
+ 8.804010000e-07 V_low
+ 8.805000000e-07 V_low
+ 8.805010000e-07 V_low
+ 8.806000000e-07 V_low
+ 8.806010000e-07 V_low
+ 8.807000000e-07 V_low
+ 8.807010000e-07 V_low
+ 8.808000000e-07 V_low
+ 8.808010000e-07 V_low
+ 8.809000000e-07 V_low
+ 8.809010000e-07 V_hig
+ 8.810000000e-07 V_hig
+ 8.810010000e-07 V_hig
+ 8.811000000e-07 V_hig
+ 8.811010000e-07 V_hig
+ 8.812000000e-07 V_hig
+ 8.812010000e-07 V_hig
+ 8.813000000e-07 V_hig
+ 8.813010000e-07 V_hig
+ 8.814000000e-07 V_hig
+ 8.814010000e-07 V_hig
+ 8.815000000e-07 V_hig
+ 8.815010000e-07 V_hig
+ 8.816000000e-07 V_hig
+ 8.816010000e-07 V_hig
+ 8.817000000e-07 V_hig
+ 8.817010000e-07 V_hig
+ 8.818000000e-07 V_hig
+ 8.818010000e-07 V_hig
+ 8.819000000e-07 V_hig
+ 8.819010000e-07 V_hig
+ 8.820000000e-07 V_hig
+ 8.820010000e-07 V_hig
+ 8.821000000e-07 V_hig
+ 8.821010000e-07 V_hig
+ 8.822000000e-07 V_hig
+ 8.822010000e-07 V_hig
+ 8.823000000e-07 V_hig
+ 8.823010000e-07 V_hig
+ 8.824000000e-07 V_hig
+ 8.824010000e-07 V_hig
+ 8.825000000e-07 V_hig
+ 8.825010000e-07 V_hig
+ 8.826000000e-07 V_hig
+ 8.826010000e-07 V_hig
+ 8.827000000e-07 V_hig
+ 8.827010000e-07 V_hig
+ 8.828000000e-07 V_hig
+ 8.828010000e-07 V_hig
+ 8.829000000e-07 V_hig
+ 8.829010000e-07 V_hig
+ 8.830000000e-07 V_hig
+ 8.830010000e-07 V_hig
+ 8.831000000e-07 V_hig
+ 8.831010000e-07 V_hig
+ 8.832000000e-07 V_hig
+ 8.832010000e-07 V_hig
+ 8.833000000e-07 V_hig
+ 8.833010000e-07 V_hig
+ 8.834000000e-07 V_hig
+ 8.834010000e-07 V_hig
+ 8.835000000e-07 V_hig
+ 8.835010000e-07 V_hig
+ 8.836000000e-07 V_hig
+ 8.836010000e-07 V_hig
+ 8.837000000e-07 V_hig
+ 8.837010000e-07 V_hig
+ 8.838000000e-07 V_hig
+ 8.838010000e-07 V_hig
+ 8.839000000e-07 V_hig
+ 8.839010000e-07 V_low
+ 8.840000000e-07 V_low
+ 8.840010000e-07 V_low
+ 8.841000000e-07 V_low
+ 8.841010000e-07 V_low
+ 8.842000000e-07 V_low
+ 8.842010000e-07 V_low
+ 8.843000000e-07 V_low
+ 8.843010000e-07 V_low
+ 8.844000000e-07 V_low
+ 8.844010000e-07 V_low
+ 8.845000000e-07 V_low
+ 8.845010000e-07 V_low
+ 8.846000000e-07 V_low
+ 8.846010000e-07 V_low
+ 8.847000000e-07 V_low
+ 8.847010000e-07 V_low
+ 8.848000000e-07 V_low
+ 8.848010000e-07 V_low
+ 8.849000000e-07 V_low
+ 8.849010000e-07 V_low
+ 8.850000000e-07 V_low
+ 8.850010000e-07 V_low
+ 8.851000000e-07 V_low
+ 8.851010000e-07 V_low
+ 8.852000000e-07 V_low
+ 8.852010000e-07 V_low
+ 8.853000000e-07 V_low
+ 8.853010000e-07 V_low
+ 8.854000000e-07 V_low
+ 8.854010000e-07 V_low
+ 8.855000000e-07 V_low
+ 8.855010000e-07 V_low
+ 8.856000000e-07 V_low
+ 8.856010000e-07 V_low
+ 8.857000000e-07 V_low
+ 8.857010000e-07 V_low
+ 8.858000000e-07 V_low
+ 8.858010000e-07 V_low
+ 8.859000000e-07 V_low
+ 8.859010000e-07 V_low
+ 8.860000000e-07 V_low
+ 8.860010000e-07 V_low
+ 8.861000000e-07 V_low
+ 8.861010000e-07 V_low
+ 8.862000000e-07 V_low
+ 8.862010000e-07 V_low
+ 8.863000000e-07 V_low
+ 8.863010000e-07 V_low
+ 8.864000000e-07 V_low
+ 8.864010000e-07 V_low
+ 8.865000000e-07 V_low
+ 8.865010000e-07 V_low
+ 8.866000000e-07 V_low
+ 8.866010000e-07 V_low
+ 8.867000000e-07 V_low
+ 8.867010000e-07 V_low
+ 8.868000000e-07 V_low
+ 8.868010000e-07 V_low
+ 8.869000000e-07 V_low
+ 8.869010000e-07 V_low
+ 8.870000000e-07 V_low
+ 8.870010000e-07 V_low
+ 8.871000000e-07 V_low
+ 8.871010000e-07 V_low
+ 8.872000000e-07 V_low
+ 8.872010000e-07 V_low
+ 8.873000000e-07 V_low
+ 8.873010000e-07 V_low
+ 8.874000000e-07 V_low
+ 8.874010000e-07 V_low
+ 8.875000000e-07 V_low
+ 8.875010000e-07 V_low
+ 8.876000000e-07 V_low
+ 8.876010000e-07 V_low
+ 8.877000000e-07 V_low
+ 8.877010000e-07 V_low
+ 8.878000000e-07 V_low
+ 8.878010000e-07 V_low
+ 8.879000000e-07 V_low
+ 8.879010000e-07 V_hig
+ 8.880000000e-07 V_hig
+ 8.880010000e-07 V_hig
+ 8.881000000e-07 V_hig
+ 8.881010000e-07 V_hig
+ 8.882000000e-07 V_hig
+ 8.882010000e-07 V_hig
+ 8.883000000e-07 V_hig
+ 8.883010000e-07 V_hig
+ 8.884000000e-07 V_hig
+ 8.884010000e-07 V_hig
+ 8.885000000e-07 V_hig
+ 8.885010000e-07 V_hig
+ 8.886000000e-07 V_hig
+ 8.886010000e-07 V_hig
+ 8.887000000e-07 V_hig
+ 8.887010000e-07 V_hig
+ 8.888000000e-07 V_hig
+ 8.888010000e-07 V_hig
+ 8.889000000e-07 V_hig
+ 8.889010000e-07 V_low
+ 8.890000000e-07 V_low
+ 8.890010000e-07 V_low
+ 8.891000000e-07 V_low
+ 8.891010000e-07 V_low
+ 8.892000000e-07 V_low
+ 8.892010000e-07 V_low
+ 8.893000000e-07 V_low
+ 8.893010000e-07 V_low
+ 8.894000000e-07 V_low
+ 8.894010000e-07 V_low
+ 8.895000000e-07 V_low
+ 8.895010000e-07 V_low
+ 8.896000000e-07 V_low
+ 8.896010000e-07 V_low
+ 8.897000000e-07 V_low
+ 8.897010000e-07 V_low
+ 8.898000000e-07 V_low
+ 8.898010000e-07 V_low
+ 8.899000000e-07 V_low
+ 8.899010000e-07 V_hig
+ 8.900000000e-07 V_hig
+ 8.900010000e-07 V_hig
+ 8.901000000e-07 V_hig
+ 8.901010000e-07 V_hig
+ 8.902000000e-07 V_hig
+ 8.902010000e-07 V_hig
+ 8.903000000e-07 V_hig
+ 8.903010000e-07 V_hig
+ 8.904000000e-07 V_hig
+ 8.904010000e-07 V_hig
+ 8.905000000e-07 V_hig
+ 8.905010000e-07 V_hig
+ 8.906000000e-07 V_hig
+ 8.906010000e-07 V_hig
+ 8.907000000e-07 V_hig
+ 8.907010000e-07 V_hig
+ 8.908000000e-07 V_hig
+ 8.908010000e-07 V_hig
+ 8.909000000e-07 V_hig
+ 8.909010000e-07 V_low
+ 8.910000000e-07 V_low
+ 8.910010000e-07 V_low
+ 8.911000000e-07 V_low
+ 8.911010000e-07 V_low
+ 8.912000000e-07 V_low
+ 8.912010000e-07 V_low
+ 8.913000000e-07 V_low
+ 8.913010000e-07 V_low
+ 8.914000000e-07 V_low
+ 8.914010000e-07 V_low
+ 8.915000000e-07 V_low
+ 8.915010000e-07 V_low
+ 8.916000000e-07 V_low
+ 8.916010000e-07 V_low
+ 8.917000000e-07 V_low
+ 8.917010000e-07 V_low
+ 8.918000000e-07 V_low
+ 8.918010000e-07 V_low
+ 8.919000000e-07 V_low
+ 8.919010000e-07 V_hig
+ 8.920000000e-07 V_hig
+ 8.920010000e-07 V_hig
+ 8.921000000e-07 V_hig
+ 8.921010000e-07 V_hig
+ 8.922000000e-07 V_hig
+ 8.922010000e-07 V_hig
+ 8.923000000e-07 V_hig
+ 8.923010000e-07 V_hig
+ 8.924000000e-07 V_hig
+ 8.924010000e-07 V_hig
+ 8.925000000e-07 V_hig
+ 8.925010000e-07 V_hig
+ 8.926000000e-07 V_hig
+ 8.926010000e-07 V_hig
+ 8.927000000e-07 V_hig
+ 8.927010000e-07 V_hig
+ 8.928000000e-07 V_hig
+ 8.928010000e-07 V_hig
+ 8.929000000e-07 V_hig
+ 8.929010000e-07 V_hig
+ 8.930000000e-07 V_hig
+ 8.930010000e-07 V_hig
+ 8.931000000e-07 V_hig
+ 8.931010000e-07 V_hig
+ 8.932000000e-07 V_hig
+ 8.932010000e-07 V_hig
+ 8.933000000e-07 V_hig
+ 8.933010000e-07 V_hig
+ 8.934000000e-07 V_hig
+ 8.934010000e-07 V_hig
+ 8.935000000e-07 V_hig
+ 8.935010000e-07 V_hig
+ 8.936000000e-07 V_hig
+ 8.936010000e-07 V_hig
+ 8.937000000e-07 V_hig
+ 8.937010000e-07 V_hig
+ 8.938000000e-07 V_hig
+ 8.938010000e-07 V_hig
+ 8.939000000e-07 V_hig
+ 8.939010000e-07 V_low
+ 8.940000000e-07 V_low
+ 8.940010000e-07 V_low
+ 8.941000000e-07 V_low
+ 8.941010000e-07 V_low
+ 8.942000000e-07 V_low
+ 8.942010000e-07 V_low
+ 8.943000000e-07 V_low
+ 8.943010000e-07 V_low
+ 8.944000000e-07 V_low
+ 8.944010000e-07 V_low
+ 8.945000000e-07 V_low
+ 8.945010000e-07 V_low
+ 8.946000000e-07 V_low
+ 8.946010000e-07 V_low
+ 8.947000000e-07 V_low
+ 8.947010000e-07 V_low
+ 8.948000000e-07 V_low
+ 8.948010000e-07 V_low
+ 8.949000000e-07 V_low
+ 8.949010000e-07 V_low
+ 8.950000000e-07 V_low
+ 8.950010000e-07 V_low
+ 8.951000000e-07 V_low
+ 8.951010000e-07 V_low
+ 8.952000000e-07 V_low
+ 8.952010000e-07 V_low
+ 8.953000000e-07 V_low
+ 8.953010000e-07 V_low
+ 8.954000000e-07 V_low
+ 8.954010000e-07 V_low
+ 8.955000000e-07 V_low
+ 8.955010000e-07 V_low
+ 8.956000000e-07 V_low
+ 8.956010000e-07 V_low
+ 8.957000000e-07 V_low
+ 8.957010000e-07 V_low
+ 8.958000000e-07 V_low
+ 8.958010000e-07 V_low
+ 8.959000000e-07 V_low
+ 8.959010000e-07 V_hig
+ 8.960000000e-07 V_hig
+ 8.960010000e-07 V_hig
+ 8.961000000e-07 V_hig
+ 8.961010000e-07 V_hig
+ 8.962000000e-07 V_hig
+ 8.962010000e-07 V_hig
+ 8.963000000e-07 V_hig
+ 8.963010000e-07 V_hig
+ 8.964000000e-07 V_hig
+ 8.964010000e-07 V_hig
+ 8.965000000e-07 V_hig
+ 8.965010000e-07 V_hig
+ 8.966000000e-07 V_hig
+ 8.966010000e-07 V_hig
+ 8.967000000e-07 V_hig
+ 8.967010000e-07 V_hig
+ 8.968000000e-07 V_hig
+ 8.968010000e-07 V_hig
+ 8.969000000e-07 V_hig
+ 8.969010000e-07 V_low
+ 8.970000000e-07 V_low
+ 8.970010000e-07 V_low
+ 8.971000000e-07 V_low
+ 8.971010000e-07 V_low
+ 8.972000000e-07 V_low
+ 8.972010000e-07 V_low
+ 8.973000000e-07 V_low
+ 8.973010000e-07 V_low
+ 8.974000000e-07 V_low
+ 8.974010000e-07 V_low
+ 8.975000000e-07 V_low
+ 8.975010000e-07 V_low
+ 8.976000000e-07 V_low
+ 8.976010000e-07 V_low
+ 8.977000000e-07 V_low
+ 8.977010000e-07 V_low
+ 8.978000000e-07 V_low
+ 8.978010000e-07 V_low
+ 8.979000000e-07 V_low
+ 8.979010000e-07 V_low
+ 8.980000000e-07 V_low
+ 8.980010000e-07 V_low
+ 8.981000000e-07 V_low
+ 8.981010000e-07 V_low
+ 8.982000000e-07 V_low
+ 8.982010000e-07 V_low
+ 8.983000000e-07 V_low
+ 8.983010000e-07 V_low
+ 8.984000000e-07 V_low
+ 8.984010000e-07 V_low
+ 8.985000000e-07 V_low
+ 8.985010000e-07 V_low
+ 8.986000000e-07 V_low
+ 8.986010000e-07 V_low
+ 8.987000000e-07 V_low
+ 8.987010000e-07 V_low
+ 8.988000000e-07 V_low
+ 8.988010000e-07 V_low
+ 8.989000000e-07 V_low
+ 8.989010000e-07 V_hig
+ 8.990000000e-07 V_hig
+ 8.990010000e-07 V_hig
+ 8.991000000e-07 V_hig
+ 8.991010000e-07 V_hig
+ 8.992000000e-07 V_hig
+ 8.992010000e-07 V_hig
+ 8.993000000e-07 V_hig
+ 8.993010000e-07 V_hig
+ 8.994000000e-07 V_hig
+ 8.994010000e-07 V_hig
+ 8.995000000e-07 V_hig
+ 8.995010000e-07 V_hig
+ 8.996000000e-07 V_hig
+ 8.996010000e-07 V_hig
+ 8.997000000e-07 V_hig
+ 8.997010000e-07 V_hig
+ 8.998000000e-07 V_hig
+ 8.998010000e-07 V_hig
+ 8.999000000e-07 V_hig
+ 8.999010000e-07 V_hig
+ 9.000000000e-07 V_hig
+ 9.000010000e-07 V_hig
+ 9.001000000e-07 V_hig
+ 9.001010000e-07 V_hig
+ 9.002000000e-07 V_hig
+ 9.002010000e-07 V_hig
+ 9.003000000e-07 V_hig
+ 9.003010000e-07 V_hig
+ 9.004000000e-07 V_hig
+ 9.004010000e-07 V_hig
+ 9.005000000e-07 V_hig
+ 9.005010000e-07 V_hig
+ 9.006000000e-07 V_hig
+ 9.006010000e-07 V_hig
+ 9.007000000e-07 V_hig
+ 9.007010000e-07 V_hig
+ 9.008000000e-07 V_hig
+ 9.008010000e-07 V_hig
+ 9.009000000e-07 V_hig
+ 9.009010000e-07 V_low
+ 9.010000000e-07 V_low
+ 9.010010000e-07 V_low
+ 9.011000000e-07 V_low
+ 9.011010000e-07 V_low
+ 9.012000000e-07 V_low
+ 9.012010000e-07 V_low
+ 9.013000000e-07 V_low
+ 9.013010000e-07 V_low
+ 9.014000000e-07 V_low
+ 9.014010000e-07 V_low
+ 9.015000000e-07 V_low
+ 9.015010000e-07 V_low
+ 9.016000000e-07 V_low
+ 9.016010000e-07 V_low
+ 9.017000000e-07 V_low
+ 9.017010000e-07 V_low
+ 9.018000000e-07 V_low
+ 9.018010000e-07 V_low
+ 9.019000000e-07 V_low
+ 9.019010000e-07 V_hig
+ 9.020000000e-07 V_hig
+ 9.020010000e-07 V_hig
+ 9.021000000e-07 V_hig
+ 9.021010000e-07 V_hig
+ 9.022000000e-07 V_hig
+ 9.022010000e-07 V_hig
+ 9.023000000e-07 V_hig
+ 9.023010000e-07 V_hig
+ 9.024000000e-07 V_hig
+ 9.024010000e-07 V_hig
+ 9.025000000e-07 V_hig
+ 9.025010000e-07 V_hig
+ 9.026000000e-07 V_hig
+ 9.026010000e-07 V_hig
+ 9.027000000e-07 V_hig
+ 9.027010000e-07 V_hig
+ 9.028000000e-07 V_hig
+ 9.028010000e-07 V_hig
+ 9.029000000e-07 V_hig
+ 9.029010000e-07 V_hig
+ 9.030000000e-07 V_hig
+ 9.030010000e-07 V_hig
+ 9.031000000e-07 V_hig
+ 9.031010000e-07 V_hig
+ 9.032000000e-07 V_hig
+ 9.032010000e-07 V_hig
+ 9.033000000e-07 V_hig
+ 9.033010000e-07 V_hig
+ 9.034000000e-07 V_hig
+ 9.034010000e-07 V_hig
+ 9.035000000e-07 V_hig
+ 9.035010000e-07 V_hig
+ 9.036000000e-07 V_hig
+ 9.036010000e-07 V_hig
+ 9.037000000e-07 V_hig
+ 9.037010000e-07 V_hig
+ 9.038000000e-07 V_hig
+ 9.038010000e-07 V_hig
+ 9.039000000e-07 V_hig
+ 9.039010000e-07 V_low
+ 9.040000000e-07 V_low
+ 9.040010000e-07 V_low
+ 9.041000000e-07 V_low
+ 9.041010000e-07 V_low
+ 9.042000000e-07 V_low
+ 9.042010000e-07 V_low
+ 9.043000000e-07 V_low
+ 9.043010000e-07 V_low
+ 9.044000000e-07 V_low
+ 9.044010000e-07 V_low
+ 9.045000000e-07 V_low
+ 9.045010000e-07 V_low
+ 9.046000000e-07 V_low
+ 9.046010000e-07 V_low
+ 9.047000000e-07 V_low
+ 9.047010000e-07 V_low
+ 9.048000000e-07 V_low
+ 9.048010000e-07 V_low
+ 9.049000000e-07 V_low
+ 9.049010000e-07 V_low
+ 9.050000000e-07 V_low
+ 9.050010000e-07 V_low
+ 9.051000000e-07 V_low
+ 9.051010000e-07 V_low
+ 9.052000000e-07 V_low
+ 9.052010000e-07 V_low
+ 9.053000000e-07 V_low
+ 9.053010000e-07 V_low
+ 9.054000000e-07 V_low
+ 9.054010000e-07 V_low
+ 9.055000000e-07 V_low
+ 9.055010000e-07 V_low
+ 9.056000000e-07 V_low
+ 9.056010000e-07 V_low
+ 9.057000000e-07 V_low
+ 9.057010000e-07 V_low
+ 9.058000000e-07 V_low
+ 9.058010000e-07 V_low
+ 9.059000000e-07 V_low
+ 9.059010000e-07 V_low
+ 9.060000000e-07 V_low
+ 9.060010000e-07 V_low
+ 9.061000000e-07 V_low
+ 9.061010000e-07 V_low
+ 9.062000000e-07 V_low
+ 9.062010000e-07 V_low
+ 9.063000000e-07 V_low
+ 9.063010000e-07 V_low
+ 9.064000000e-07 V_low
+ 9.064010000e-07 V_low
+ 9.065000000e-07 V_low
+ 9.065010000e-07 V_low
+ 9.066000000e-07 V_low
+ 9.066010000e-07 V_low
+ 9.067000000e-07 V_low
+ 9.067010000e-07 V_low
+ 9.068000000e-07 V_low
+ 9.068010000e-07 V_low
+ 9.069000000e-07 V_low
+ 9.069010000e-07 V_low
+ 9.070000000e-07 V_low
+ 9.070010000e-07 V_low
+ 9.071000000e-07 V_low
+ 9.071010000e-07 V_low
+ 9.072000000e-07 V_low
+ 9.072010000e-07 V_low
+ 9.073000000e-07 V_low
+ 9.073010000e-07 V_low
+ 9.074000000e-07 V_low
+ 9.074010000e-07 V_low
+ 9.075000000e-07 V_low
+ 9.075010000e-07 V_low
+ 9.076000000e-07 V_low
+ 9.076010000e-07 V_low
+ 9.077000000e-07 V_low
+ 9.077010000e-07 V_low
+ 9.078000000e-07 V_low
+ 9.078010000e-07 V_low
+ 9.079000000e-07 V_low
+ 9.079010000e-07 V_hig
+ 9.080000000e-07 V_hig
+ 9.080010000e-07 V_hig
+ 9.081000000e-07 V_hig
+ 9.081010000e-07 V_hig
+ 9.082000000e-07 V_hig
+ 9.082010000e-07 V_hig
+ 9.083000000e-07 V_hig
+ 9.083010000e-07 V_hig
+ 9.084000000e-07 V_hig
+ 9.084010000e-07 V_hig
+ 9.085000000e-07 V_hig
+ 9.085010000e-07 V_hig
+ 9.086000000e-07 V_hig
+ 9.086010000e-07 V_hig
+ 9.087000000e-07 V_hig
+ 9.087010000e-07 V_hig
+ 9.088000000e-07 V_hig
+ 9.088010000e-07 V_hig
+ 9.089000000e-07 V_hig
+ 9.089010000e-07 V_low
+ 9.090000000e-07 V_low
+ 9.090010000e-07 V_low
+ 9.091000000e-07 V_low
+ 9.091010000e-07 V_low
+ 9.092000000e-07 V_low
+ 9.092010000e-07 V_low
+ 9.093000000e-07 V_low
+ 9.093010000e-07 V_low
+ 9.094000000e-07 V_low
+ 9.094010000e-07 V_low
+ 9.095000000e-07 V_low
+ 9.095010000e-07 V_low
+ 9.096000000e-07 V_low
+ 9.096010000e-07 V_low
+ 9.097000000e-07 V_low
+ 9.097010000e-07 V_low
+ 9.098000000e-07 V_low
+ 9.098010000e-07 V_low
+ 9.099000000e-07 V_low
+ 9.099010000e-07 V_low
+ 9.100000000e-07 V_low
+ 9.100010000e-07 V_low
+ 9.101000000e-07 V_low
+ 9.101010000e-07 V_low
+ 9.102000000e-07 V_low
+ 9.102010000e-07 V_low
+ 9.103000000e-07 V_low
+ 9.103010000e-07 V_low
+ 9.104000000e-07 V_low
+ 9.104010000e-07 V_low
+ 9.105000000e-07 V_low
+ 9.105010000e-07 V_low
+ 9.106000000e-07 V_low
+ 9.106010000e-07 V_low
+ 9.107000000e-07 V_low
+ 9.107010000e-07 V_low
+ 9.108000000e-07 V_low
+ 9.108010000e-07 V_low
+ 9.109000000e-07 V_low
+ 9.109010000e-07 V_low
+ 9.110000000e-07 V_low
+ 9.110010000e-07 V_low
+ 9.111000000e-07 V_low
+ 9.111010000e-07 V_low
+ 9.112000000e-07 V_low
+ 9.112010000e-07 V_low
+ 9.113000000e-07 V_low
+ 9.113010000e-07 V_low
+ 9.114000000e-07 V_low
+ 9.114010000e-07 V_low
+ 9.115000000e-07 V_low
+ 9.115010000e-07 V_low
+ 9.116000000e-07 V_low
+ 9.116010000e-07 V_low
+ 9.117000000e-07 V_low
+ 9.117010000e-07 V_low
+ 9.118000000e-07 V_low
+ 9.118010000e-07 V_low
+ 9.119000000e-07 V_low
+ 9.119010000e-07 V_hig
+ 9.120000000e-07 V_hig
+ 9.120010000e-07 V_hig
+ 9.121000000e-07 V_hig
+ 9.121010000e-07 V_hig
+ 9.122000000e-07 V_hig
+ 9.122010000e-07 V_hig
+ 9.123000000e-07 V_hig
+ 9.123010000e-07 V_hig
+ 9.124000000e-07 V_hig
+ 9.124010000e-07 V_hig
+ 9.125000000e-07 V_hig
+ 9.125010000e-07 V_hig
+ 9.126000000e-07 V_hig
+ 9.126010000e-07 V_hig
+ 9.127000000e-07 V_hig
+ 9.127010000e-07 V_hig
+ 9.128000000e-07 V_hig
+ 9.128010000e-07 V_hig
+ 9.129000000e-07 V_hig
+ 9.129010000e-07 V_low
+ 9.130000000e-07 V_low
+ 9.130010000e-07 V_low
+ 9.131000000e-07 V_low
+ 9.131010000e-07 V_low
+ 9.132000000e-07 V_low
+ 9.132010000e-07 V_low
+ 9.133000000e-07 V_low
+ 9.133010000e-07 V_low
+ 9.134000000e-07 V_low
+ 9.134010000e-07 V_low
+ 9.135000000e-07 V_low
+ 9.135010000e-07 V_low
+ 9.136000000e-07 V_low
+ 9.136010000e-07 V_low
+ 9.137000000e-07 V_low
+ 9.137010000e-07 V_low
+ 9.138000000e-07 V_low
+ 9.138010000e-07 V_low
+ 9.139000000e-07 V_low
+ 9.139010000e-07 V_low
+ 9.140000000e-07 V_low
+ 9.140010000e-07 V_low
+ 9.141000000e-07 V_low
+ 9.141010000e-07 V_low
+ 9.142000000e-07 V_low
+ 9.142010000e-07 V_low
+ 9.143000000e-07 V_low
+ 9.143010000e-07 V_low
+ 9.144000000e-07 V_low
+ 9.144010000e-07 V_low
+ 9.145000000e-07 V_low
+ 9.145010000e-07 V_low
+ 9.146000000e-07 V_low
+ 9.146010000e-07 V_low
+ 9.147000000e-07 V_low
+ 9.147010000e-07 V_low
+ 9.148000000e-07 V_low
+ 9.148010000e-07 V_low
+ 9.149000000e-07 V_low
+ 9.149010000e-07 V_hig
+ 9.150000000e-07 V_hig
+ 9.150010000e-07 V_hig
+ 9.151000000e-07 V_hig
+ 9.151010000e-07 V_hig
+ 9.152000000e-07 V_hig
+ 9.152010000e-07 V_hig
+ 9.153000000e-07 V_hig
+ 9.153010000e-07 V_hig
+ 9.154000000e-07 V_hig
+ 9.154010000e-07 V_hig
+ 9.155000000e-07 V_hig
+ 9.155010000e-07 V_hig
+ 9.156000000e-07 V_hig
+ 9.156010000e-07 V_hig
+ 9.157000000e-07 V_hig
+ 9.157010000e-07 V_hig
+ 9.158000000e-07 V_hig
+ 9.158010000e-07 V_hig
+ 9.159000000e-07 V_hig
+ 9.159010000e-07 V_low
+ 9.160000000e-07 V_low
+ 9.160010000e-07 V_low
+ 9.161000000e-07 V_low
+ 9.161010000e-07 V_low
+ 9.162000000e-07 V_low
+ 9.162010000e-07 V_low
+ 9.163000000e-07 V_low
+ 9.163010000e-07 V_low
+ 9.164000000e-07 V_low
+ 9.164010000e-07 V_low
+ 9.165000000e-07 V_low
+ 9.165010000e-07 V_low
+ 9.166000000e-07 V_low
+ 9.166010000e-07 V_low
+ 9.167000000e-07 V_low
+ 9.167010000e-07 V_low
+ 9.168000000e-07 V_low
+ 9.168010000e-07 V_low
+ 9.169000000e-07 V_low
+ 9.169010000e-07 V_hig
+ 9.170000000e-07 V_hig
+ 9.170010000e-07 V_hig
+ 9.171000000e-07 V_hig
+ 9.171010000e-07 V_hig
+ 9.172000000e-07 V_hig
+ 9.172010000e-07 V_hig
+ 9.173000000e-07 V_hig
+ 9.173010000e-07 V_hig
+ 9.174000000e-07 V_hig
+ 9.174010000e-07 V_hig
+ 9.175000000e-07 V_hig
+ 9.175010000e-07 V_hig
+ 9.176000000e-07 V_hig
+ 9.176010000e-07 V_hig
+ 9.177000000e-07 V_hig
+ 9.177010000e-07 V_hig
+ 9.178000000e-07 V_hig
+ 9.178010000e-07 V_hig
+ 9.179000000e-07 V_hig
+ 9.179010000e-07 V_hig
+ 9.180000000e-07 V_hig
+ 9.180010000e-07 V_hig
+ 9.181000000e-07 V_hig
+ 9.181010000e-07 V_hig
+ 9.182000000e-07 V_hig
+ 9.182010000e-07 V_hig
+ 9.183000000e-07 V_hig
+ 9.183010000e-07 V_hig
+ 9.184000000e-07 V_hig
+ 9.184010000e-07 V_hig
+ 9.185000000e-07 V_hig
+ 9.185010000e-07 V_hig
+ 9.186000000e-07 V_hig
+ 9.186010000e-07 V_hig
+ 9.187000000e-07 V_hig
+ 9.187010000e-07 V_hig
+ 9.188000000e-07 V_hig
+ 9.188010000e-07 V_hig
+ 9.189000000e-07 V_hig
+ 9.189010000e-07 V_hig
+ 9.190000000e-07 V_hig
+ 9.190010000e-07 V_hig
+ 9.191000000e-07 V_hig
+ 9.191010000e-07 V_hig
+ 9.192000000e-07 V_hig
+ 9.192010000e-07 V_hig
+ 9.193000000e-07 V_hig
+ 9.193010000e-07 V_hig
+ 9.194000000e-07 V_hig
+ 9.194010000e-07 V_hig
+ 9.195000000e-07 V_hig
+ 9.195010000e-07 V_hig
+ 9.196000000e-07 V_hig
+ 9.196010000e-07 V_hig
+ 9.197000000e-07 V_hig
+ 9.197010000e-07 V_hig
+ 9.198000000e-07 V_hig
+ 9.198010000e-07 V_hig
+ 9.199000000e-07 V_hig
+ 9.199010000e-07 V_hig
+ 9.200000000e-07 V_hig
+ 9.200010000e-07 V_hig
+ 9.201000000e-07 V_hig
+ 9.201010000e-07 V_hig
+ 9.202000000e-07 V_hig
+ 9.202010000e-07 V_hig
+ 9.203000000e-07 V_hig
+ 9.203010000e-07 V_hig
+ 9.204000000e-07 V_hig
+ 9.204010000e-07 V_hig
+ 9.205000000e-07 V_hig
+ 9.205010000e-07 V_hig
+ 9.206000000e-07 V_hig
+ 9.206010000e-07 V_hig
+ 9.207000000e-07 V_hig
+ 9.207010000e-07 V_hig
+ 9.208000000e-07 V_hig
+ 9.208010000e-07 V_hig
+ 9.209000000e-07 V_hig
+ 9.209010000e-07 V_low
+ 9.210000000e-07 V_low
+ 9.210010000e-07 V_low
+ 9.211000000e-07 V_low
+ 9.211010000e-07 V_low
+ 9.212000000e-07 V_low
+ 9.212010000e-07 V_low
+ 9.213000000e-07 V_low
+ 9.213010000e-07 V_low
+ 9.214000000e-07 V_low
+ 9.214010000e-07 V_low
+ 9.215000000e-07 V_low
+ 9.215010000e-07 V_low
+ 9.216000000e-07 V_low
+ 9.216010000e-07 V_low
+ 9.217000000e-07 V_low
+ 9.217010000e-07 V_low
+ 9.218000000e-07 V_low
+ 9.218010000e-07 V_low
+ 9.219000000e-07 V_low
+ 9.219010000e-07 V_low
+ 9.220000000e-07 V_low
+ 9.220010000e-07 V_low
+ 9.221000000e-07 V_low
+ 9.221010000e-07 V_low
+ 9.222000000e-07 V_low
+ 9.222010000e-07 V_low
+ 9.223000000e-07 V_low
+ 9.223010000e-07 V_low
+ 9.224000000e-07 V_low
+ 9.224010000e-07 V_low
+ 9.225000000e-07 V_low
+ 9.225010000e-07 V_low
+ 9.226000000e-07 V_low
+ 9.226010000e-07 V_low
+ 9.227000000e-07 V_low
+ 9.227010000e-07 V_low
+ 9.228000000e-07 V_low
+ 9.228010000e-07 V_low
+ 9.229000000e-07 V_low
+ 9.229010000e-07 V_hig
+ 9.230000000e-07 V_hig
+ 9.230010000e-07 V_hig
+ 9.231000000e-07 V_hig
+ 9.231010000e-07 V_hig
+ 9.232000000e-07 V_hig
+ 9.232010000e-07 V_hig
+ 9.233000000e-07 V_hig
+ 9.233010000e-07 V_hig
+ 9.234000000e-07 V_hig
+ 9.234010000e-07 V_hig
+ 9.235000000e-07 V_hig
+ 9.235010000e-07 V_hig
+ 9.236000000e-07 V_hig
+ 9.236010000e-07 V_hig
+ 9.237000000e-07 V_hig
+ 9.237010000e-07 V_hig
+ 9.238000000e-07 V_hig
+ 9.238010000e-07 V_hig
+ 9.239000000e-07 V_hig
+ 9.239010000e-07 V_hig
+ 9.240000000e-07 V_hig
+ 9.240010000e-07 V_hig
+ 9.241000000e-07 V_hig
+ 9.241010000e-07 V_hig
+ 9.242000000e-07 V_hig
+ 9.242010000e-07 V_hig
+ 9.243000000e-07 V_hig
+ 9.243010000e-07 V_hig
+ 9.244000000e-07 V_hig
+ 9.244010000e-07 V_hig
+ 9.245000000e-07 V_hig
+ 9.245010000e-07 V_hig
+ 9.246000000e-07 V_hig
+ 9.246010000e-07 V_hig
+ 9.247000000e-07 V_hig
+ 9.247010000e-07 V_hig
+ 9.248000000e-07 V_hig
+ 9.248010000e-07 V_hig
+ 9.249000000e-07 V_hig
+ 9.249010000e-07 V_low
+ 9.250000000e-07 V_low
+ 9.250010000e-07 V_low
+ 9.251000000e-07 V_low
+ 9.251010000e-07 V_low
+ 9.252000000e-07 V_low
+ 9.252010000e-07 V_low
+ 9.253000000e-07 V_low
+ 9.253010000e-07 V_low
+ 9.254000000e-07 V_low
+ 9.254010000e-07 V_low
+ 9.255000000e-07 V_low
+ 9.255010000e-07 V_low
+ 9.256000000e-07 V_low
+ 9.256010000e-07 V_low
+ 9.257000000e-07 V_low
+ 9.257010000e-07 V_low
+ 9.258000000e-07 V_low
+ 9.258010000e-07 V_low
+ 9.259000000e-07 V_low
+ 9.259010000e-07 V_low
+ 9.260000000e-07 V_low
+ 9.260010000e-07 V_low
+ 9.261000000e-07 V_low
+ 9.261010000e-07 V_low
+ 9.262000000e-07 V_low
+ 9.262010000e-07 V_low
+ 9.263000000e-07 V_low
+ 9.263010000e-07 V_low
+ 9.264000000e-07 V_low
+ 9.264010000e-07 V_low
+ 9.265000000e-07 V_low
+ 9.265010000e-07 V_low
+ 9.266000000e-07 V_low
+ 9.266010000e-07 V_low
+ 9.267000000e-07 V_low
+ 9.267010000e-07 V_low
+ 9.268000000e-07 V_low
+ 9.268010000e-07 V_low
+ 9.269000000e-07 V_low
+ 9.269010000e-07 V_hig
+ 9.270000000e-07 V_hig
+ 9.270010000e-07 V_hig
+ 9.271000000e-07 V_hig
+ 9.271010000e-07 V_hig
+ 9.272000000e-07 V_hig
+ 9.272010000e-07 V_hig
+ 9.273000000e-07 V_hig
+ 9.273010000e-07 V_hig
+ 9.274000000e-07 V_hig
+ 9.274010000e-07 V_hig
+ 9.275000000e-07 V_hig
+ 9.275010000e-07 V_hig
+ 9.276000000e-07 V_hig
+ 9.276010000e-07 V_hig
+ 9.277000000e-07 V_hig
+ 9.277010000e-07 V_hig
+ 9.278000000e-07 V_hig
+ 9.278010000e-07 V_hig
+ 9.279000000e-07 V_hig
+ 9.279010000e-07 V_hig
+ 9.280000000e-07 V_hig
+ 9.280010000e-07 V_hig
+ 9.281000000e-07 V_hig
+ 9.281010000e-07 V_hig
+ 9.282000000e-07 V_hig
+ 9.282010000e-07 V_hig
+ 9.283000000e-07 V_hig
+ 9.283010000e-07 V_hig
+ 9.284000000e-07 V_hig
+ 9.284010000e-07 V_hig
+ 9.285000000e-07 V_hig
+ 9.285010000e-07 V_hig
+ 9.286000000e-07 V_hig
+ 9.286010000e-07 V_hig
+ 9.287000000e-07 V_hig
+ 9.287010000e-07 V_hig
+ 9.288000000e-07 V_hig
+ 9.288010000e-07 V_hig
+ 9.289000000e-07 V_hig
+ 9.289010000e-07 V_hig
+ 9.290000000e-07 V_hig
+ 9.290010000e-07 V_hig
+ 9.291000000e-07 V_hig
+ 9.291010000e-07 V_hig
+ 9.292000000e-07 V_hig
+ 9.292010000e-07 V_hig
+ 9.293000000e-07 V_hig
+ 9.293010000e-07 V_hig
+ 9.294000000e-07 V_hig
+ 9.294010000e-07 V_hig
+ 9.295000000e-07 V_hig
+ 9.295010000e-07 V_hig
+ 9.296000000e-07 V_hig
+ 9.296010000e-07 V_hig
+ 9.297000000e-07 V_hig
+ 9.297010000e-07 V_hig
+ 9.298000000e-07 V_hig
+ 9.298010000e-07 V_hig
+ 9.299000000e-07 V_hig
+ 9.299010000e-07 V_hig
+ 9.300000000e-07 V_hig
+ 9.300010000e-07 V_hig
+ 9.301000000e-07 V_hig
+ 9.301010000e-07 V_hig
+ 9.302000000e-07 V_hig
+ 9.302010000e-07 V_hig
+ 9.303000000e-07 V_hig
+ 9.303010000e-07 V_hig
+ 9.304000000e-07 V_hig
+ 9.304010000e-07 V_hig
+ 9.305000000e-07 V_hig
+ 9.305010000e-07 V_hig
+ 9.306000000e-07 V_hig
+ 9.306010000e-07 V_hig
+ 9.307000000e-07 V_hig
+ 9.307010000e-07 V_hig
+ 9.308000000e-07 V_hig
+ 9.308010000e-07 V_hig
+ 9.309000000e-07 V_hig
+ 9.309010000e-07 V_hig
+ 9.310000000e-07 V_hig
+ 9.310010000e-07 V_hig
+ 9.311000000e-07 V_hig
+ 9.311010000e-07 V_hig
+ 9.312000000e-07 V_hig
+ 9.312010000e-07 V_hig
+ 9.313000000e-07 V_hig
+ 9.313010000e-07 V_hig
+ 9.314000000e-07 V_hig
+ 9.314010000e-07 V_hig
+ 9.315000000e-07 V_hig
+ 9.315010000e-07 V_hig
+ 9.316000000e-07 V_hig
+ 9.316010000e-07 V_hig
+ 9.317000000e-07 V_hig
+ 9.317010000e-07 V_hig
+ 9.318000000e-07 V_hig
+ 9.318010000e-07 V_hig
+ 9.319000000e-07 V_hig
+ 9.319010000e-07 V_low
+ 9.320000000e-07 V_low
+ 9.320010000e-07 V_low
+ 9.321000000e-07 V_low
+ 9.321010000e-07 V_low
+ 9.322000000e-07 V_low
+ 9.322010000e-07 V_low
+ 9.323000000e-07 V_low
+ 9.323010000e-07 V_low
+ 9.324000000e-07 V_low
+ 9.324010000e-07 V_low
+ 9.325000000e-07 V_low
+ 9.325010000e-07 V_low
+ 9.326000000e-07 V_low
+ 9.326010000e-07 V_low
+ 9.327000000e-07 V_low
+ 9.327010000e-07 V_low
+ 9.328000000e-07 V_low
+ 9.328010000e-07 V_low
+ 9.329000000e-07 V_low
+ 9.329010000e-07 V_hig
+ 9.330000000e-07 V_hig
+ 9.330010000e-07 V_hig
+ 9.331000000e-07 V_hig
+ 9.331010000e-07 V_hig
+ 9.332000000e-07 V_hig
+ 9.332010000e-07 V_hig
+ 9.333000000e-07 V_hig
+ 9.333010000e-07 V_hig
+ 9.334000000e-07 V_hig
+ 9.334010000e-07 V_hig
+ 9.335000000e-07 V_hig
+ 9.335010000e-07 V_hig
+ 9.336000000e-07 V_hig
+ 9.336010000e-07 V_hig
+ 9.337000000e-07 V_hig
+ 9.337010000e-07 V_hig
+ 9.338000000e-07 V_hig
+ 9.338010000e-07 V_hig
+ 9.339000000e-07 V_hig
+ 9.339010000e-07 V_low
+ 9.340000000e-07 V_low
+ 9.340010000e-07 V_low
+ 9.341000000e-07 V_low
+ 9.341010000e-07 V_low
+ 9.342000000e-07 V_low
+ 9.342010000e-07 V_low
+ 9.343000000e-07 V_low
+ 9.343010000e-07 V_low
+ 9.344000000e-07 V_low
+ 9.344010000e-07 V_low
+ 9.345000000e-07 V_low
+ 9.345010000e-07 V_low
+ 9.346000000e-07 V_low
+ 9.346010000e-07 V_low
+ 9.347000000e-07 V_low
+ 9.347010000e-07 V_low
+ 9.348000000e-07 V_low
+ 9.348010000e-07 V_low
+ 9.349000000e-07 V_low
+ 9.349010000e-07 V_hig
+ 9.350000000e-07 V_hig
+ 9.350010000e-07 V_hig
+ 9.351000000e-07 V_hig
+ 9.351010000e-07 V_hig
+ 9.352000000e-07 V_hig
+ 9.352010000e-07 V_hig
+ 9.353000000e-07 V_hig
+ 9.353010000e-07 V_hig
+ 9.354000000e-07 V_hig
+ 9.354010000e-07 V_hig
+ 9.355000000e-07 V_hig
+ 9.355010000e-07 V_hig
+ 9.356000000e-07 V_hig
+ 9.356010000e-07 V_hig
+ 9.357000000e-07 V_hig
+ 9.357010000e-07 V_hig
+ 9.358000000e-07 V_hig
+ 9.358010000e-07 V_hig
+ 9.359000000e-07 V_hig
+ 9.359010000e-07 V_low
+ 9.360000000e-07 V_low
+ 9.360010000e-07 V_low
+ 9.361000000e-07 V_low
+ 9.361010000e-07 V_low
+ 9.362000000e-07 V_low
+ 9.362010000e-07 V_low
+ 9.363000000e-07 V_low
+ 9.363010000e-07 V_low
+ 9.364000000e-07 V_low
+ 9.364010000e-07 V_low
+ 9.365000000e-07 V_low
+ 9.365010000e-07 V_low
+ 9.366000000e-07 V_low
+ 9.366010000e-07 V_low
+ 9.367000000e-07 V_low
+ 9.367010000e-07 V_low
+ 9.368000000e-07 V_low
+ 9.368010000e-07 V_low
+ 9.369000000e-07 V_low
+ 9.369010000e-07 V_low
+ 9.370000000e-07 V_low
+ 9.370010000e-07 V_low
+ 9.371000000e-07 V_low
+ 9.371010000e-07 V_low
+ 9.372000000e-07 V_low
+ 9.372010000e-07 V_low
+ 9.373000000e-07 V_low
+ 9.373010000e-07 V_low
+ 9.374000000e-07 V_low
+ 9.374010000e-07 V_low
+ 9.375000000e-07 V_low
+ 9.375010000e-07 V_low
+ 9.376000000e-07 V_low
+ 9.376010000e-07 V_low
+ 9.377000000e-07 V_low
+ 9.377010000e-07 V_low
+ 9.378000000e-07 V_low
+ 9.378010000e-07 V_low
+ 9.379000000e-07 V_low
+ 9.379010000e-07 V_hig
+ 9.380000000e-07 V_hig
+ 9.380010000e-07 V_hig
+ 9.381000000e-07 V_hig
+ 9.381010000e-07 V_hig
+ 9.382000000e-07 V_hig
+ 9.382010000e-07 V_hig
+ 9.383000000e-07 V_hig
+ 9.383010000e-07 V_hig
+ 9.384000000e-07 V_hig
+ 9.384010000e-07 V_hig
+ 9.385000000e-07 V_hig
+ 9.385010000e-07 V_hig
+ 9.386000000e-07 V_hig
+ 9.386010000e-07 V_hig
+ 9.387000000e-07 V_hig
+ 9.387010000e-07 V_hig
+ 9.388000000e-07 V_hig
+ 9.388010000e-07 V_hig
+ 9.389000000e-07 V_hig
+ 9.389010000e-07 V_hig
+ 9.390000000e-07 V_hig
+ 9.390010000e-07 V_hig
+ 9.391000000e-07 V_hig
+ 9.391010000e-07 V_hig
+ 9.392000000e-07 V_hig
+ 9.392010000e-07 V_hig
+ 9.393000000e-07 V_hig
+ 9.393010000e-07 V_hig
+ 9.394000000e-07 V_hig
+ 9.394010000e-07 V_hig
+ 9.395000000e-07 V_hig
+ 9.395010000e-07 V_hig
+ 9.396000000e-07 V_hig
+ 9.396010000e-07 V_hig
+ 9.397000000e-07 V_hig
+ 9.397010000e-07 V_hig
+ 9.398000000e-07 V_hig
+ 9.398010000e-07 V_hig
+ 9.399000000e-07 V_hig
+ 9.399010000e-07 V_hig
+ 9.400000000e-07 V_hig
+ 9.400010000e-07 V_hig
+ 9.401000000e-07 V_hig
+ 9.401010000e-07 V_hig
+ 9.402000000e-07 V_hig
+ 9.402010000e-07 V_hig
+ 9.403000000e-07 V_hig
+ 9.403010000e-07 V_hig
+ 9.404000000e-07 V_hig
+ 9.404010000e-07 V_hig
+ 9.405000000e-07 V_hig
+ 9.405010000e-07 V_hig
+ 9.406000000e-07 V_hig
+ 9.406010000e-07 V_hig
+ 9.407000000e-07 V_hig
+ 9.407010000e-07 V_hig
+ 9.408000000e-07 V_hig
+ 9.408010000e-07 V_hig
+ 9.409000000e-07 V_hig
+ 9.409010000e-07 V_low
+ 9.410000000e-07 V_low
+ 9.410010000e-07 V_low
+ 9.411000000e-07 V_low
+ 9.411010000e-07 V_low
+ 9.412000000e-07 V_low
+ 9.412010000e-07 V_low
+ 9.413000000e-07 V_low
+ 9.413010000e-07 V_low
+ 9.414000000e-07 V_low
+ 9.414010000e-07 V_low
+ 9.415000000e-07 V_low
+ 9.415010000e-07 V_low
+ 9.416000000e-07 V_low
+ 9.416010000e-07 V_low
+ 9.417000000e-07 V_low
+ 9.417010000e-07 V_low
+ 9.418000000e-07 V_low
+ 9.418010000e-07 V_low
+ 9.419000000e-07 V_low
+ 9.419010000e-07 V_low
+ 9.420000000e-07 V_low
+ 9.420010000e-07 V_low
+ 9.421000000e-07 V_low
+ 9.421010000e-07 V_low
+ 9.422000000e-07 V_low
+ 9.422010000e-07 V_low
+ 9.423000000e-07 V_low
+ 9.423010000e-07 V_low
+ 9.424000000e-07 V_low
+ 9.424010000e-07 V_low
+ 9.425000000e-07 V_low
+ 9.425010000e-07 V_low
+ 9.426000000e-07 V_low
+ 9.426010000e-07 V_low
+ 9.427000000e-07 V_low
+ 9.427010000e-07 V_low
+ 9.428000000e-07 V_low
+ 9.428010000e-07 V_low
+ 9.429000000e-07 V_low
+ 9.429010000e-07 V_hig
+ 9.430000000e-07 V_hig
+ 9.430010000e-07 V_hig
+ 9.431000000e-07 V_hig
+ 9.431010000e-07 V_hig
+ 9.432000000e-07 V_hig
+ 9.432010000e-07 V_hig
+ 9.433000000e-07 V_hig
+ 9.433010000e-07 V_hig
+ 9.434000000e-07 V_hig
+ 9.434010000e-07 V_hig
+ 9.435000000e-07 V_hig
+ 9.435010000e-07 V_hig
+ 9.436000000e-07 V_hig
+ 9.436010000e-07 V_hig
+ 9.437000000e-07 V_hig
+ 9.437010000e-07 V_hig
+ 9.438000000e-07 V_hig
+ 9.438010000e-07 V_hig
+ 9.439000000e-07 V_hig
+ 9.439010000e-07 V_hig
+ 9.440000000e-07 V_hig
+ 9.440010000e-07 V_hig
+ 9.441000000e-07 V_hig
+ 9.441010000e-07 V_hig
+ 9.442000000e-07 V_hig
+ 9.442010000e-07 V_hig
+ 9.443000000e-07 V_hig
+ 9.443010000e-07 V_hig
+ 9.444000000e-07 V_hig
+ 9.444010000e-07 V_hig
+ 9.445000000e-07 V_hig
+ 9.445010000e-07 V_hig
+ 9.446000000e-07 V_hig
+ 9.446010000e-07 V_hig
+ 9.447000000e-07 V_hig
+ 9.447010000e-07 V_hig
+ 9.448000000e-07 V_hig
+ 9.448010000e-07 V_hig
+ 9.449000000e-07 V_hig
+ 9.449010000e-07 V_low
+ 9.450000000e-07 V_low
+ 9.450010000e-07 V_low
+ 9.451000000e-07 V_low
+ 9.451010000e-07 V_low
+ 9.452000000e-07 V_low
+ 9.452010000e-07 V_low
+ 9.453000000e-07 V_low
+ 9.453010000e-07 V_low
+ 9.454000000e-07 V_low
+ 9.454010000e-07 V_low
+ 9.455000000e-07 V_low
+ 9.455010000e-07 V_low
+ 9.456000000e-07 V_low
+ 9.456010000e-07 V_low
+ 9.457000000e-07 V_low
+ 9.457010000e-07 V_low
+ 9.458000000e-07 V_low
+ 9.458010000e-07 V_low
+ 9.459000000e-07 V_low
+ 9.459010000e-07 V_low
+ 9.460000000e-07 V_low
+ 9.460010000e-07 V_low
+ 9.461000000e-07 V_low
+ 9.461010000e-07 V_low
+ 9.462000000e-07 V_low
+ 9.462010000e-07 V_low
+ 9.463000000e-07 V_low
+ 9.463010000e-07 V_low
+ 9.464000000e-07 V_low
+ 9.464010000e-07 V_low
+ 9.465000000e-07 V_low
+ 9.465010000e-07 V_low
+ 9.466000000e-07 V_low
+ 9.466010000e-07 V_low
+ 9.467000000e-07 V_low
+ 9.467010000e-07 V_low
+ 9.468000000e-07 V_low
+ 9.468010000e-07 V_low
+ 9.469000000e-07 V_low
+ 9.469010000e-07 V_low
+ 9.470000000e-07 V_low
+ 9.470010000e-07 V_low
+ 9.471000000e-07 V_low
+ 9.471010000e-07 V_low
+ 9.472000000e-07 V_low
+ 9.472010000e-07 V_low
+ 9.473000000e-07 V_low
+ 9.473010000e-07 V_low
+ 9.474000000e-07 V_low
+ 9.474010000e-07 V_low
+ 9.475000000e-07 V_low
+ 9.475010000e-07 V_low
+ 9.476000000e-07 V_low
+ 9.476010000e-07 V_low
+ 9.477000000e-07 V_low
+ 9.477010000e-07 V_low
+ 9.478000000e-07 V_low
+ 9.478010000e-07 V_low
+ 9.479000000e-07 V_low
+ 9.479010000e-07 V_low
+ 9.480000000e-07 V_low
+ 9.480010000e-07 V_low
+ 9.481000000e-07 V_low
+ 9.481010000e-07 V_low
+ 9.482000000e-07 V_low
+ 9.482010000e-07 V_low
+ 9.483000000e-07 V_low
+ 9.483010000e-07 V_low
+ 9.484000000e-07 V_low
+ 9.484010000e-07 V_low
+ 9.485000000e-07 V_low
+ 9.485010000e-07 V_low
+ 9.486000000e-07 V_low
+ 9.486010000e-07 V_low
+ 9.487000000e-07 V_low
+ 9.487010000e-07 V_low
+ 9.488000000e-07 V_low
+ 9.488010000e-07 V_low
+ 9.489000000e-07 V_low
+ 9.489010000e-07 V_hig
+ 9.490000000e-07 V_hig
+ 9.490010000e-07 V_hig
+ 9.491000000e-07 V_hig
+ 9.491010000e-07 V_hig
+ 9.492000000e-07 V_hig
+ 9.492010000e-07 V_hig
+ 9.493000000e-07 V_hig
+ 9.493010000e-07 V_hig
+ 9.494000000e-07 V_hig
+ 9.494010000e-07 V_hig
+ 9.495000000e-07 V_hig
+ 9.495010000e-07 V_hig
+ 9.496000000e-07 V_hig
+ 9.496010000e-07 V_hig
+ 9.497000000e-07 V_hig
+ 9.497010000e-07 V_hig
+ 9.498000000e-07 V_hig
+ 9.498010000e-07 V_hig
+ 9.499000000e-07 V_hig
+ 9.499010000e-07 V_hig
+ 9.500000000e-07 V_hig
+ 9.500010000e-07 V_hig
+ 9.501000000e-07 V_hig
+ 9.501010000e-07 V_hig
+ 9.502000000e-07 V_hig
+ 9.502010000e-07 V_hig
+ 9.503000000e-07 V_hig
+ 9.503010000e-07 V_hig
+ 9.504000000e-07 V_hig
+ 9.504010000e-07 V_hig
+ 9.505000000e-07 V_hig
+ 9.505010000e-07 V_hig
+ 9.506000000e-07 V_hig
+ 9.506010000e-07 V_hig
+ 9.507000000e-07 V_hig
+ 9.507010000e-07 V_hig
+ 9.508000000e-07 V_hig
+ 9.508010000e-07 V_hig
+ 9.509000000e-07 V_hig
+ 9.509010000e-07 V_low
+ 9.510000000e-07 V_low
+ 9.510010000e-07 V_low
+ 9.511000000e-07 V_low
+ 9.511010000e-07 V_low
+ 9.512000000e-07 V_low
+ 9.512010000e-07 V_low
+ 9.513000000e-07 V_low
+ 9.513010000e-07 V_low
+ 9.514000000e-07 V_low
+ 9.514010000e-07 V_low
+ 9.515000000e-07 V_low
+ 9.515010000e-07 V_low
+ 9.516000000e-07 V_low
+ 9.516010000e-07 V_low
+ 9.517000000e-07 V_low
+ 9.517010000e-07 V_low
+ 9.518000000e-07 V_low
+ 9.518010000e-07 V_low
+ 9.519000000e-07 V_low
+ 9.519010000e-07 V_hig
+ 9.520000000e-07 V_hig
+ 9.520010000e-07 V_hig
+ 9.521000000e-07 V_hig
+ 9.521010000e-07 V_hig
+ 9.522000000e-07 V_hig
+ 9.522010000e-07 V_hig
+ 9.523000000e-07 V_hig
+ 9.523010000e-07 V_hig
+ 9.524000000e-07 V_hig
+ 9.524010000e-07 V_hig
+ 9.525000000e-07 V_hig
+ 9.525010000e-07 V_hig
+ 9.526000000e-07 V_hig
+ 9.526010000e-07 V_hig
+ 9.527000000e-07 V_hig
+ 9.527010000e-07 V_hig
+ 9.528000000e-07 V_hig
+ 9.528010000e-07 V_hig
+ 9.529000000e-07 V_hig
+ 9.529010000e-07 V_low
+ 9.530000000e-07 V_low
+ 9.530010000e-07 V_low
+ 9.531000000e-07 V_low
+ 9.531010000e-07 V_low
+ 9.532000000e-07 V_low
+ 9.532010000e-07 V_low
+ 9.533000000e-07 V_low
+ 9.533010000e-07 V_low
+ 9.534000000e-07 V_low
+ 9.534010000e-07 V_low
+ 9.535000000e-07 V_low
+ 9.535010000e-07 V_low
+ 9.536000000e-07 V_low
+ 9.536010000e-07 V_low
+ 9.537000000e-07 V_low
+ 9.537010000e-07 V_low
+ 9.538000000e-07 V_low
+ 9.538010000e-07 V_low
+ 9.539000000e-07 V_low
+ 9.539010000e-07 V_low
+ 9.540000000e-07 V_low
+ 9.540010000e-07 V_low
+ 9.541000000e-07 V_low
+ 9.541010000e-07 V_low
+ 9.542000000e-07 V_low
+ 9.542010000e-07 V_low
+ 9.543000000e-07 V_low
+ 9.543010000e-07 V_low
+ 9.544000000e-07 V_low
+ 9.544010000e-07 V_low
+ 9.545000000e-07 V_low
+ 9.545010000e-07 V_low
+ 9.546000000e-07 V_low
+ 9.546010000e-07 V_low
+ 9.547000000e-07 V_low
+ 9.547010000e-07 V_low
+ 9.548000000e-07 V_low
+ 9.548010000e-07 V_low
+ 9.549000000e-07 V_low
+ 9.549010000e-07 V_hig
+ 9.550000000e-07 V_hig
+ 9.550010000e-07 V_hig
+ 9.551000000e-07 V_hig
+ 9.551010000e-07 V_hig
+ 9.552000000e-07 V_hig
+ 9.552010000e-07 V_hig
+ 9.553000000e-07 V_hig
+ 9.553010000e-07 V_hig
+ 9.554000000e-07 V_hig
+ 9.554010000e-07 V_hig
+ 9.555000000e-07 V_hig
+ 9.555010000e-07 V_hig
+ 9.556000000e-07 V_hig
+ 9.556010000e-07 V_hig
+ 9.557000000e-07 V_hig
+ 9.557010000e-07 V_hig
+ 9.558000000e-07 V_hig
+ 9.558010000e-07 V_hig
+ 9.559000000e-07 V_hig
+ 9.559010000e-07 V_hig
+ 9.560000000e-07 V_hig
+ 9.560010000e-07 V_hig
+ 9.561000000e-07 V_hig
+ 9.561010000e-07 V_hig
+ 9.562000000e-07 V_hig
+ 9.562010000e-07 V_hig
+ 9.563000000e-07 V_hig
+ 9.563010000e-07 V_hig
+ 9.564000000e-07 V_hig
+ 9.564010000e-07 V_hig
+ 9.565000000e-07 V_hig
+ 9.565010000e-07 V_hig
+ 9.566000000e-07 V_hig
+ 9.566010000e-07 V_hig
+ 9.567000000e-07 V_hig
+ 9.567010000e-07 V_hig
+ 9.568000000e-07 V_hig
+ 9.568010000e-07 V_hig
+ 9.569000000e-07 V_hig
+ 9.569010000e-07 V_low
+ 9.570000000e-07 V_low
+ 9.570010000e-07 V_low
+ 9.571000000e-07 V_low
+ 9.571010000e-07 V_low
+ 9.572000000e-07 V_low
+ 9.572010000e-07 V_low
+ 9.573000000e-07 V_low
+ 9.573010000e-07 V_low
+ 9.574000000e-07 V_low
+ 9.574010000e-07 V_low
+ 9.575000000e-07 V_low
+ 9.575010000e-07 V_low
+ 9.576000000e-07 V_low
+ 9.576010000e-07 V_low
+ 9.577000000e-07 V_low
+ 9.577010000e-07 V_low
+ 9.578000000e-07 V_low
+ 9.578010000e-07 V_low
+ 9.579000000e-07 V_low
+ 9.579010000e-07 V_low
+ 9.580000000e-07 V_low
+ 9.580010000e-07 V_low
+ 9.581000000e-07 V_low
+ 9.581010000e-07 V_low
+ 9.582000000e-07 V_low
+ 9.582010000e-07 V_low
+ 9.583000000e-07 V_low
+ 9.583010000e-07 V_low
+ 9.584000000e-07 V_low
+ 9.584010000e-07 V_low
+ 9.585000000e-07 V_low
+ 9.585010000e-07 V_low
+ 9.586000000e-07 V_low
+ 9.586010000e-07 V_low
+ 9.587000000e-07 V_low
+ 9.587010000e-07 V_low
+ 9.588000000e-07 V_low
+ 9.588010000e-07 V_low
+ 9.589000000e-07 V_low
+ 9.589010000e-07 V_low
+ 9.590000000e-07 V_low
+ 9.590010000e-07 V_low
+ 9.591000000e-07 V_low
+ 9.591010000e-07 V_low
+ 9.592000000e-07 V_low
+ 9.592010000e-07 V_low
+ 9.593000000e-07 V_low
+ 9.593010000e-07 V_low
+ 9.594000000e-07 V_low
+ 9.594010000e-07 V_low
+ 9.595000000e-07 V_low
+ 9.595010000e-07 V_low
+ 9.596000000e-07 V_low
+ 9.596010000e-07 V_low
+ 9.597000000e-07 V_low
+ 9.597010000e-07 V_low
+ 9.598000000e-07 V_low
+ 9.598010000e-07 V_low
+ 9.599000000e-07 V_low
+ 9.599010000e-07 V_low
+ 9.600000000e-07 V_low
+ 9.600010000e-07 V_low
+ 9.601000000e-07 V_low
+ 9.601010000e-07 V_low
+ 9.602000000e-07 V_low
+ 9.602010000e-07 V_low
+ 9.603000000e-07 V_low
+ 9.603010000e-07 V_low
+ 9.604000000e-07 V_low
+ 9.604010000e-07 V_low
+ 9.605000000e-07 V_low
+ 9.605010000e-07 V_low
+ 9.606000000e-07 V_low
+ 9.606010000e-07 V_low
+ 9.607000000e-07 V_low
+ 9.607010000e-07 V_low
+ 9.608000000e-07 V_low
+ 9.608010000e-07 V_low
+ 9.609000000e-07 V_low
+ 9.609010000e-07 V_low
+ 9.610000000e-07 V_low
+ 9.610010000e-07 V_low
+ 9.611000000e-07 V_low
+ 9.611010000e-07 V_low
+ 9.612000000e-07 V_low
+ 9.612010000e-07 V_low
+ 9.613000000e-07 V_low
+ 9.613010000e-07 V_low
+ 9.614000000e-07 V_low
+ 9.614010000e-07 V_low
+ 9.615000000e-07 V_low
+ 9.615010000e-07 V_low
+ 9.616000000e-07 V_low
+ 9.616010000e-07 V_low
+ 9.617000000e-07 V_low
+ 9.617010000e-07 V_low
+ 9.618000000e-07 V_low
+ 9.618010000e-07 V_low
+ 9.619000000e-07 V_low
+ 9.619010000e-07 V_hig
+ 9.620000000e-07 V_hig
+ 9.620010000e-07 V_hig
+ 9.621000000e-07 V_hig
+ 9.621010000e-07 V_hig
+ 9.622000000e-07 V_hig
+ 9.622010000e-07 V_hig
+ 9.623000000e-07 V_hig
+ 9.623010000e-07 V_hig
+ 9.624000000e-07 V_hig
+ 9.624010000e-07 V_hig
+ 9.625000000e-07 V_hig
+ 9.625010000e-07 V_hig
+ 9.626000000e-07 V_hig
+ 9.626010000e-07 V_hig
+ 9.627000000e-07 V_hig
+ 9.627010000e-07 V_hig
+ 9.628000000e-07 V_hig
+ 9.628010000e-07 V_hig
+ 9.629000000e-07 V_hig
+ 9.629010000e-07 V_hig
+ 9.630000000e-07 V_hig
+ 9.630010000e-07 V_hig
+ 9.631000000e-07 V_hig
+ 9.631010000e-07 V_hig
+ 9.632000000e-07 V_hig
+ 9.632010000e-07 V_hig
+ 9.633000000e-07 V_hig
+ 9.633010000e-07 V_hig
+ 9.634000000e-07 V_hig
+ 9.634010000e-07 V_hig
+ 9.635000000e-07 V_hig
+ 9.635010000e-07 V_hig
+ 9.636000000e-07 V_hig
+ 9.636010000e-07 V_hig
+ 9.637000000e-07 V_hig
+ 9.637010000e-07 V_hig
+ 9.638000000e-07 V_hig
+ 9.638010000e-07 V_hig
+ 9.639000000e-07 V_hig
+ 9.639010000e-07 V_low
+ 9.640000000e-07 V_low
+ 9.640010000e-07 V_low
+ 9.641000000e-07 V_low
+ 9.641010000e-07 V_low
+ 9.642000000e-07 V_low
+ 9.642010000e-07 V_low
+ 9.643000000e-07 V_low
+ 9.643010000e-07 V_low
+ 9.644000000e-07 V_low
+ 9.644010000e-07 V_low
+ 9.645000000e-07 V_low
+ 9.645010000e-07 V_low
+ 9.646000000e-07 V_low
+ 9.646010000e-07 V_low
+ 9.647000000e-07 V_low
+ 9.647010000e-07 V_low
+ 9.648000000e-07 V_low
+ 9.648010000e-07 V_low
+ 9.649000000e-07 V_low
+ 9.649010000e-07 V_low
+ 9.650000000e-07 V_low
+ 9.650010000e-07 V_low
+ 9.651000000e-07 V_low
+ 9.651010000e-07 V_low
+ 9.652000000e-07 V_low
+ 9.652010000e-07 V_low
+ 9.653000000e-07 V_low
+ 9.653010000e-07 V_low
+ 9.654000000e-07 V_low
+ 9.654010000e-07 V_low
+ 9.655000000e-07 V_low
+ 9.655010000e-07 V_low
+ 9.656000000e-07 V_low
+ 9.656010000e-07 V_low
+ 9.657000000e-07 V_low
+ 9.657010000e-07 V_low
+ 9.658000000e-07 V_low
+ 9.658010000e-07 V_low
+ 9.659000000e-07 V_low
+ 9.659010000e-07 V_hig
+ 9.660000000e-07 V_hig
+ 9.660010000e-07 V_hig
+ 9.661000000e-07 V_hig
+ 9.661010000e-07 V_hig
+ 9.662000000e-07 V_hig
+ 9.662010000e-07 V_hig
+ 9.663000000e-07 V_hig
+ 9.663010000e-07 V_hig
+ 9.664000000e-07 V_hig
+ 9.664010000e-07 V_hig
+ 9.665000000e-07 V_hig
+ 9.665010000e-07 V_hig
+ 9.666000000e-07 V_hig
+ 9.666010000e-07 V_hig
+ 9.667000000e-07 V_hig
+ 9.667010000e-07 V_hig
+ 9.668000000e-07 V_hig
+ 9.668010000e-07 V_hig
+ 9.669000000e-07 V_hig
+ 9.669010000e-07 V_low
+ 9.670000000e-07 V_low
+ 9.670010000e-07 V_low
+ 9.671000000e-07 V_low
+ 9.671010000e-07 V_low
+ 9.672000000e-07 V_low
+ 9.672010000e-07 V_low
+ 9.673000000e-07 V_low
+ 9.673010000e-07 V_low
+ 9.674000000e-07 V_low
+ 9.674010000e-07 V_low
+ 9.675000000e-07 V_low
+ 9.675010000e-07 V_low
+ 9.676000000e-07 V_low
+ 9.676010000e-07 V_low
+ 9.677000000e-07 V_low
+ 9.677010000e-07 V_low
+ 9.678000000e-07 V_low
+ 9.678010000e-07 V_low
+ 9.679000000e-07 V_low
+ 9.679010000e-07 V_hig
+ 9.680000000e-07 V_hig
+ 9.680010000e-07 V_hig
+ 9.681000000e-07 V_hig
+ 9.681010000e-07 V_hig
+ 9.682000000e-07 V_hig
+ 9.682010000e-07 V_hig
+ 9.683000000e-07 V_hig
+ 9.683010000e-07 V_hig
+ 9.684000000e-07 V_hig
+ 9.684010000e-07 V_hig
+ 9.685000000e-07 V_hig
+ 9.685010000e-07 V_hig
+ 9.686000000e-07 V_hig
+ 9.686010000e-07 V_hig
+ 9.687000000e-07 V_hig
+ 9.687010000e-07 V_hig
+ 9.688000000e-07 V_hig
+ 9.688010000e-07 V_hig
+ 9.689000000e-07 V_hig
+ 9.689010000e-07 V_hig
+ 9.690000000e-07 V_hig
+ 9.690010000e-07 V_hig
+ 9.691000000e-07 V_hig
+ 9.691010000e-07 V_hig
+ 9.692000000e-07 V_hig
+ 9.692010000e-07 V_hig
+ 9.693000000e-07 V_hig
+ 9.693010000e-07 V_hig
+ 9.694000000e-07 V_hig
+ 9.694010000e-07 V_hig
+ 9.695000000e-07 V_hig
+ 9.695010000e-07 V_hig
+ 9.696000000e-07 V_hig
+ 9.696010000e-07 V_hig
+ 9.697000000e-07 V_hig
+ 9.697010000e-07 V_hig
+ 9.698000000e-07 V_hig
+ 9.698010000e-07 V_hig
+ 9.699000000e-07 V_hig
+ 9.699010000e-07 V_low
+ 9.700000000e-07 V_low
+ 9.700010000e-07 V_low
+ 9.701000000e-07 V_low
+ 9.701010000e-07 V_low
+ 9.702000000e-07 V_low
+ 9.702010000e-07 V_low
+ 9.703000000e-07 V_low
+ 9.703010000e-07 V_low
+ 9.704000000e-07 V_low
+ 9.704010000e-07 V_low
+ 9.705000000e-07 V_low
+ 9.705010000e-07 V_low
+ 9.706000000e-07 V_low
+ 9.706010000e-07 V_low
+ 9.707000000e-07 V_low
+ 9.707010000e-07 V_low
+ 9.708000000e-07 V_low
+ 9.708010000e-07 V_low
+ 9.709000000e-07 V_low
+ 9.709010000e-07 V_low
+ 9.710000000e-07 V_low
+ 9.710010000e-07 V_low
+ 9.711000000e-07 V_low
+ 9.711010000e-07 V_low
+ 9.712000000e-07 V_low
+ 9.712010000e-07 V_low
+ 9.713000000e-07 V_low
+ 9.713010000e-07 V_low
+ 9.714000000e-07 V_low
+ 9.714010000e-07 V_low
+ 9.715000000e-07 V_low
+ 9.715010000e-07 V_low
+ 9.716000000e-07 V_low
+ 9.716010000e-07 V_low
+ 9.717000000e-07 V_low
+ 9.717010000e-07 V_low
+ 9.718000000e-07 V_low
+ 9.718010000e-07 V_low
+ 9.719000000e-07 V_low
+ 9.719010000e-07 V_hig
+ 9.720000000e-07 V_hig
+ 9.720010000e-07 V_hig
+ 9.721000000e-07 V_hig
+ 9.721010000e-07 V_hig
+ 9.722000000e-07 V_hig
+ 9.722010000e-07 V_hig
+ 9.723000000e-07 V_hig
+ 9.723010000e-07 V_hig
+ 9.724000000e-07 V_hig
+ 9.724010000e-07 V_hig
+ 9.725000000e-07 V_hig
+ 9.725010000e-07 V_hig
+ 9.726000000e-07 V_hig
+ 9.726010000e-07 V_hig
+ 9.727000000e-07 V_hig
+ 9.727010000e-07 V_hig
+ 9.728000000e-07 V_hig
+ 9.728010000e-07 V_hig
+ 9.729000000e-07 V_hig
+ 9.729010000e-07 V_low
+ 9.730000000e-07 V_low
+ 9.730010000e-07 V_low
+ 9.731000000e-07 V_low
+ 9.731010000e-07 V_low
+ 9.732000000e-07 V_low
+ 9.732010000e-07 V_low
+ 9.733000000e-07 V_low
+ 9.733010000e-07 V_low
+ 9.734000000e-07 V_low
+ 9.734010000e-07 V_low
+ 9.735000000e-07 V_low
+ 9.735010000e-07 V_low
+ 9.736000000e-07 V_low
+ 9.736010000e-07 V_low
+ 9.737000000e-07 V_low
+ 9.737010000e-07 V_low
+ 9.738000000e-07 V_low
+ 9.738010000e-07 V_low
+ 9.739000000e-07 V_low
+ 9.739010000e-07 V_low
+ 9.740000000e-07 V_low
+ 9.740010000e-07 V_low
+ 9.741000000e-07 V_low
+ 9.741010000e-07 V_low
+ 9.742000000e-07 V_low
+ 9.742010000e-07 V_low
+ 9.743000000e-07 V_low
+ 9.743010000e-07 V_low
+ 9.744000000e-07 V_low
+ 9.744010000e-07 V_low
+ 9.745000000e-07 V_low
+ 9.745010000e-07 V_low
+ 9.746000000e-07 V_low
+ 9.746010000e-07 V_low
+ 9.747000000e-07 V_low
+ 9.747010000e-07 V_low
+ 9.748000000e-07 V_low
+ 9.748010000e-07 V_low
+ 9.749000000e-07 V_low
+ 9.749010000e-07 V_low
+ 9.750000000e-07 V_low
+ 9.750010000e-07 V_low
+ 9.751000000e-07 V_low
+ 9.751010000e-07 V_low
+ 9.752000000e-07 V_low
+ 9.752010000e-07 V_low
+ 9.753000000e-07 V_low
+ 9.753010000e-07 V_low
+ 9.754000000e-07 V_low
+ 9.754010000e-07 V_low
+ 9.755000000e-07 V_low
+ 9.755010000e-07 V_low
+ 9.756000000e-07 V_low
+ 9.756010000e-07 V_low
+ 9.757000000e-07 V_low
+ 9.757010000e-07 V_low
+ 9.758000000e-07 V_low
+ 9.758010000e-07 V_low
+ 9.759000000e-07 V_low
+ 9.759010000e-07 V_hig
+ 9.760000000e-07 V_hig
+ 9.760010000e-07 V_hig
+ 9.761000000e-07 V_hig
+ 9.761010000e-07 V_hig
+ 9.762000000e-07 V_hig
+ 9.762010000e-07 V_hig
+ 9.763000000e-07 V_hig
+ 9.763010000e-07 V_hig
+ 9.764000000e-07 V_hig
+ 9.764010000e-07 V_hig
+ 9.765000000e-07 V_hig
+ 9.765010000e-07 V_hig
+ 9.766000000e-07 V_hig
+ 9.766010000e-07 V_hig
+ 9.767000000e-07 V_hig
+ 9.767010000e-07 V_hig
+ 9.768000000e-07 V_hig
+ 9.768010000e-07 V_hig
+ 9.769000000e-07 V_hig
+ 9.769010000e-07 V_hig
+ 9.770000000e-07 V_hig
+ 9.770010000e-07 V_hig
+ 9.771000000e-07 V_hig
+ 9.771010000e-07 V_hig
+ 9.772000000e-07 V_hig
+ 9.772010000e-07 V_hig
+ 9.773000000e-07 V_hig
+ 9.773010000e-07 V_hig
+ 9.774000000e-07 V_hig
+ 9.774010000e-07 V_hig
+ 9.775000000e-07 V_hig
+ 9.775010000e-07 V_hig
+ 9.776000000e-07 V_hig
+ 9.776010000e-07 V_hig
+ 9.777000000e-07 V_hig
+ 9.777010000e-07 V_hig
+ 9.778000000e-07 V_hig
+ 9.778010000e-07 V_hig
+ 9.779000000e-07 V_hig
+ 9.779010000e-07 V_low
+ 9.780000000e-07 V_low
+ 9.780010000e-07 V_low
+ 9.781000000e-07 V_low
+ 9.781010000e-07 V_low
+ 9.782000000e-07 V_low
+ 9.782010000e-07 V_low
+ 9.783000000e-07 V_low
+ 9.783010000e-07 V_low
+ 9.784000000e-07 V_low
+ 9.784010000e-07 V_low
+ 9.785000000e-07 V_low
+ 9.785010000e-07 V_low
+ 9.786000000e-07 V_low
+ 9.786010000e-07 V_low
+ 9.787000000e-07 V_low
+ 9.787010000e-07 V_low
+ 9.788000000e-07 V_low
+ 9.788010000e-07 V_low
+ 9.789000000e-07 V_low
+ 9.789010000e-07 V_hig
+ 9.790000000e-07 V_hig
+ 9.790010000e-07 V_hig
+ 9.791000000e-07 V_hig
+ 9.791010000e-07 V_hig
+ 9.792000000e-07 V_hig
+ 9.792010000e-07 V_hig
+ 9.793000000e-07 V_hig
+ 9.793010000e-07 V_hig
+ 9.794000000e-07 V_hig
+ 9.794010000e-07 V_hig
+ 9.795000000e-07 V_hig
+ 9.795010000e-07 V_hig
+ 9.796000000e-07 V_hig
+ 9.796010000e-07 V_hig
+ 9.797000000e-07 V_hig
+ 9.797010000e-07 V_hig
+ 9.798000000e-07 V_hig
+ 9.798010000e-07 V_hig
+ 9.799000000e-07 V_hig
+ 9.799010000e-07 V_hig
+ 9.800000000e-07 V_hig
+ 9.800010000e-07 V_hig
+ 9.801000000e-07 V_hig
+ 9.801010000e-07 V_hig
+ 9.802000000e-07 V_hig
+ 9.802010000e-07 V_hig
+ 9.803000000e-07 V_hig
+ 9.803010000e-07 V_hig
+ 9.804000000e-07 V_hig
+ 9.804010000e-07 V_hig
+ 9.805000000e-07 V_hig
+ 9.805010000e-07 V_hig
+ 9.806000000e-07 V_hig
+ 9.806010000e-07 V_hig
+ 9.807000000e-07 V_hig
+ 9.807010000e-07 V_hig
+ 9.808000000e-07 V_hig
+ 9.808010000e-07 V_hig
+ 9.809000000e-07 V_hig
+ 9.809010000e-07 V_hig
+ 9.810000000e-07 V_hig
+ 9.810010000e-07 V_hig
+ 9.811000000e-07 V_hig
+ 9.811010000e-07 V_hig
+ 9.812000000e-07 V_hig
+ 9.812010000e-07 V_hig
+ 9.813000000e-07 V_hig
+ 9.813010000e-07 V_hig
+ 9.814000000e-07 V_hig
+ 9.814010000e-07 V_hig
+ 9.815000000e-07 V_hig
+ 9.815010000e-07 V_hig
+ 9.816000000e-07 V_hig
+ 9.816010000e-07 V_hig
+ 9.817000000e-07 V_hig
+ 9.817010000e-07 V_hig
+ 9.818000000e-07 V_hig
+ 9.818010000e-07 V_hig
+ 9.819000000e-07 V_hig
+ 9.819010000e-07 V_low
+ 9.820000000e-07 V_low
+ 9.820010000e-07 V_low
+ 9.821000000e-07 V_low
+ 9.821010000e-07 V_low
+ 9.822000000e-07 V_low
+ 9.822010000e-07 V_low
+ 9.823000000e-07 V_low
+ 9.823010000e-07 V_low
+ 9.824000000e-07 V_low
+ 9.824010000e-07 V_low
+ 9.825000000e-07 V_low
+ 9.825010000e-07 V_low
+ 9.826000000e-07 V_low
+ 9.826010000e-07 V_low
+ 9.827000000e-07 V_low
+ 9.827010000e-07 V_low
+ 9.828000000e-07 V_low
+ 9.828010000e-07 V_low
+ 9.829000000e-07 V_low
+ 9.829010000e-07 V_hig
+ 9.830000000e-07 V_hig
+ 9.830010000e-07 V_hig
+ 9.831000000e-07 V_hig
+ 9.831010000e-07 V_hig
+ 9.832000000e-07 V_hig
+ 9.832010000e-07 V_hig
+ 9.833000000e-07 V_hig
+ 9.833010000e-07 V_hig
+ 9.834000000e-07 V_hig
+ 9.834010000e-07 V_hig
+ 9.835000000e-07 V_hig
+ 9.835010000e-07 V_hig
+ 9.836000000e-07 V_hig
+ 9.836010000e-07 V_hig
+ 9.837000000e-07 V_hig
+ 9.837010000e-07 V_hig
+ 9.838000000e-07 V_hig
+ 9.838010000e-07 V_hig
+ 9.839000000e-07 V_hig
+ 9.839010000e-07 V_low
+ 9.840000000e-07 V_low
+ 9.840010000e-07 V_low
+ 9.841000000e-07 V_low
+ 9.841010000e-07 V_low
+ 9.842000000e-07 V_low
+ 9.842010000e-07 V_low
+ 9.843000000e-07 V_low
+ 9.843010000e-07 V_low
+ 9.844000000e-07 V_low
+ 9.844010000e-07 V_low
+ 9.845000000e-07 V_low
+ 9.845010000e-07 V_low
+ 9.846000000e-07 V_low
+ 9.846010000e-07 V_low
+ 9.847000000e-07 V_low
+ 9.847010000e-07 V_low
+ 9.848000000e-07 V_low
+ 9.848010000e-07 V_low
+ 9.849000000e-07 V_low
+ 9.849010000e-07 V_hig
+ 9.850000000e-07 V_hig
+ 9.850010000e-07 V_hig
+ 9.851000000e-07 V_hig
+ 9.851010000e-07 V_hig
+ 9.852000000e-07 V_hig
+ 9.852010000e-07 V_hig
+ 9.853000000e-07 V_hig
+ 9.853010000e-07 V_hig
+ 9.854000000e-07 V_hig
+ 9.854010000e-07 V_hig
+ 9.855000000e-07 V_hig
+ 9.855010000e-07 V_hig
+ 9.856000000e-07 V_hig
+ 9.856010000e-07 V_hig
+ 9.857000000e-07 V_hig
+ 9.857010000e-07 V_hig
+ 9.858000000e-07 V_hig
+ 9.858010000e-07 V_hig
+ 9.859000000e-07 V_hig
+ 9.859010000e-07 V_hig
+ 9.860000000e-07 V_hig
+ 9.860010000e-07 V_hig
+ 9.861000000e-07 V_hig
+ 9.861010000e-07 V_hig
+ 9.862000000e-07 V_hig
+ 9.862010000e-07 V_hig
+ 9.863000000e-07 V_hig
+ 9.863010000e-07 V_hig
+ 9.864000000e-07 V_hig
+ 9.864010000e-07 V_hig
+ 9.865000000e-07 V_hig
+ 9.865010000e-07 V_hig
+ 9.866000000e-07 V_hig
+ 9.866010000e-07 V_hig
+ 9.867000000e-07 V_hig
+ 9.867010000e-07 V_hig
+ 9.868000000e-07 V_hig
+ 9.868010000e-07 V_hig
+ 9.869000000e-07 V_hig
+ 9.869010000e-07 V_low
+ 9.870000000e-07 V_low
+ 9.870010000e-07 V_low
+ 9.871000000e-07 V_low
+ 9.871010000e-07 V_low
+ 9.872000000e-07 V_low
+ 9.872010000e-07 V_low
+ 9.873000000e-07 V_low
+ 9.873010000e-07 V_low
+ 9.874000000e-07 V_low
+ 9.874010000e-07 V_low
+ 9.875000000e-07 V_low
+ 9.875010000e-07 V_low
+ 9.876000000e-07 V_low
+ 9.876010000e-07 V_low
+ 9.877000000e-07 V_low
+ 9.877010000e-07 V_low
+ 9.878000000e-07 V_low
+ 9.878010000e-07 V_low
+ 9.879000000e-07 V_low
+ 9.879010000e-07 V_low
+ 9.880000000e-07 V_low
+ 9.880010000e-07 V_low
+ 9.881000000e-07 V_low
+ 9.881010000e-07 V_low
+ 9.882000000e-07 V_low
+ 9.882010000e-07 V_low
+ 9.883000000e-07 V_low
+ 9.883010000e-07 V_low
+ 9.884000000e-07 V_low
+ 9.884010000e-07 V_low
+ 9.885000000e-07 V_low
+ 9.885010000e-07 V_low
+ 9.886000000e-07 V_low
+ 9.886010000e-07 V_low
+ 9.887000000e-07 V_low
+ 9.887010000e-07 V_low
+ 9.888000000e-07 V_low
+ 9.888010000e-07 V_low
+ 9.889000000e-07 V_low
+ 9.889010000e-07 V_low
+ 9.890000000e-07 V_low
+ 9.890010000e-07 V_low
+ 9.891000000e-07 V_low
+ 9.891010000e-07 V_low
+ 9.892000000e-07 V_low
+ 9.892010000e-07 V_low
+ 9.893000000e-07 V_low
+ 9.893010000e-07 V_low
+ 9.894000000e-07 V_low
+ 9.894010000e-07 V_low
+ 9.895000000e-07 V_low
+ 9.895010000e-07 V_low
+ 9.896000000e-07 V_low
+ 9.896010000e-07 V_low
+ 9.897000000e-07 V_low
+ 9.897010000e-07 V_low
+ 9.898000000e-07 V_low
+ 9.898010000e-07 V_low
+ 9.899000000e-07 V_low
+ 9.899010000e-07 V_low
+ 9.900000000e-07 V_low
+ 9.900010000e-07 V_low
+ 9.901000000e-07 V_low
+ 9.901010000e-07 V_low
+ 9.902000000e-07 V_low
+ 9.902010000e-07 V_low
+ 9.903000000e-07 V_low
+ 9.903010000e-07 V_low
+ 9.904000000e-07 V_low
+ 9.904010000e-07 V_low
+ 9.905000000e-07 V_low
+ 9.905010000e-07 V_low
+ 9.906000000e-07 V_low
+ 9.906010000e-07 V_low
+ 9.907000000e-07 V_low
+ 9.907010000e-07 V_low
+ 9.908000000e-07 V_low
+ 9.908010000e-07 V_low
+ 9.909000000e-07 V_low
+ 9.909010000e-07 V_hig
+ 9.910000000e-07 V_hig
+ 9.910010000e-07 V_hig
+ 9.911000000e-07 V_hig
+ 9.911010000e-07 V_hig
+ 9.912000000e-07 V_hig
+ 9.912010000e-07 V_hig
+ 9.913000000e-07 V_hig
+ 9.913010000e-07 V_hig
+ 9.914000000e-07 V_hig
+ 9.914010000e-07 V_hig
+ 9.915000000e-07 V_hig
+ 9.915010000e-07 V_hig
+ 9.916000000e-07 V_hig
+ 9.916010000e-07 V_hig
+ 9.917000000e-07 V_hig
+ 9.917010000e-07 V_hig
+ 9.918000000e-07 V_hig
+ 9.918010000e-07 V_hig
+ 9.919000000e-07 V_hig
+ 9.919010000e-07 V_hig
+ 9.920000000e-07 V_hig
+ 9.920010000e-07 V_hig
+ 9.921000000e-07 V_hig
+ 9.921010000e-07 V_hig
+ 9.922000000e-07 V_hig
+ 9.922010000e-07 V_hig
+ 9.923000000e-07 V_hig
+ 9.923010000e-07 V_hig
+ 9.924000000e-07 V_hig
+ 9.924010000e-07 V_hig
+ 9.925000000e-07 V_hig
+ 9.925010000e-07 V_hig
+ 9.926000000e-07 V_hig
+ 9.926010000e-07 V_hig
+ 9.927000000e-07 V_hig
+ 9.927010000e-07 V_hig
+ 9.928000000e-07 V_hig
+ 9.928010000e-07 V_hig
+ 9.929000000e-07 V_hig
+ 9.929010000e-07 V_hig
+ 9.930000000e-07 V_hig
+ 9.930010000e-07 V_hig
+ 9.931000000e-07 V_hig
+ 9.931010000e-07 V_hig
+ 9.932000000e-07 V_hig
+ 9.932010000e-07 V_hig
+ 9.933000000e-07 V_hig
+ 9.933010000e-07 V_hig
+ 9.934000000e-07 V_hig
+ 9.934010000e-07 V_hig
+ 9.935000000e-07 V_hig
+ 9.935010000e-07 V_hig
+ 9.936000000e-07 V_hig
+ 9.936010000e-07 V_hig
+ 9.937000000e-07 V_hig
+ 9.937010000e-07 V_hig
+ 9.938000000e-07 V_hig
+ 9.938010000e-07 V_hig
+ 9.939000000e-07 V_hig
+ 9.939010000e-07 V_low
+ 9.940000000e-07 V_low
+ 9.940010000e-07 V_low
+ 9.941000000e-07 V_low
+ 9.941010000e-07 V_low
+ 9.942000000e-07 V_low
+ 9.942010000e-07 V_low
+ 9.943000000e-07 V_low
+ 9.943010000e-07 V_low
+ 9.944000000e-07 V_low
+ 9.944010000e-07 V_low
+ 9.945000000e-07 V_low
+ 9.945010000e-07 V_low
+ 9.946000000e-07 V_low
+ 9.946010000e-07 V_low
+ 9.947000000e-07 V_low
+ 9.947010000e-07 V_low
+ 9.948000000e-07 V_low
+ 9.948010000e-07 V_low
+ 9.949000000e-07 V_low
+ 9.949010000e-07 V_hig
+ 9.950000000e-07 V_hig
+ 9.950010000e-07 V_hig
+ 9.951000000e-07 V_hig
+ 9.951010000e-07 V_hig
+ 9.952000000e-07 V_hig
+ 9.952010000e-07 V_hig
+ 9.953000000e-07 V_hig
+ 9.953010000e-07 V_hig
+ 9.954000000e-07 V_hig
+ 9.954010000e-07 V_hig
+ 9.955000000e-07 V_hig
+ 9.955010000e-07 V_hig
+ 9.956000000e-07 V_hig
+ 9.956010000e-07 V_hig
+ 9.957000000e-07 V_hig
+ 9.957010000e-07 V_hig
+ 9.958000000e-07 V_hig
+ 9.958010000e-07 V_hig
+ 9.959000000e-07 V_hig
+ 9.959010000e-07 V_hig
+ 9.960000000e-07 V_hig
+ 9.960010000e-07 V_hig
+ 9.961000000e-07 V_hig
+ 9.961010000e-07 V_hig
+ 9.962000000e-07 V_hig
+ 9.962010000e-07 V_hig
+ 9.963000000e-07 V_hig
+ 9.963010000e-07 V_hig
+ 9.964000000e-07 V_hig
+ 9.964010000e-07 V_hig
+ 9.965000000e-07 V_hig
+ 9.965010000e-07 V_hig
+ 9.966000000e-07 V_hig
+ 9.966010000e-07 V_hig
+ 9.967000000e-07 V_hig
+ 9.967010000e-07 V_hig
+ 9.968000000e-07 V_hig
+ 9.968010000e-07 V_hig
+ 9.969000000e-07 V_hig
+ 9.969010000e-07 V_hig
+ 9.970000000e-07 V_hig
+ 9.970010000e-07 V_hig
+ 9.971000000e-07 V_hig
+ 9.971010000e-07 V_hig
+ 9.972000000e-07 V_hig
+ 9.972010000e-07 V_hig
+ 9.973000000e-07 V_hig
+ 9.973010000e-07 V_hig
+ 9.974000000e-07 V_hig
+ 9.974010000e-07 V_hig
+ 9.975000000e-07 V_hig
+ 9.975010000e-07 V_hig
+ 9.976000000e-07 V_hig
+ 9.976010000e-07 V_hig
+ 9.977000000e-07 V_hig
+ 9.977010000e-07 V_hig
+ 9.978000000e-07 V_hig
+ 9.978010000e-07 V_hig
+ 9.979000000e-07 V_hig
+ 9.979010000e-07 V_hig
+ 9.980000000e-07 V_hig
+ 9.980010000e-07 V_hig
+ 9.981000000e-07 V_hig
+ 9.981010000e-07 V_hig
+ 9.982000000e-07 V_hig
+ 9.982010000e-07 V_hig
+ 9.983000000e-07 V_hig
+ 9.983010000e-07 V_hig
+ 9.984000000e-07 V_hig
+ 9.984010000e-07 V_hig
+ 9.985000000e-07 V_hig
+ 9.985010000e-07 V_hig
+ 9.986000000e-07 V_hig
+ 9.986010000e-07 V_hig
+ 9.987000000e-07 V_hig
+ 9.987010000e-07 V_hig
+ 9.988000000e-07 V_hig
+ 9.988010000e-07 V_hig
+ 9.989000000e-07 V_hig
+ 9.989010000e-07 V_low
+ 9.990000000e-07 V_low
+ 9.990010000e-07 V_low
+ 9.991000000e-07 V_low
+ 9.991010000e-07 V_low
+ 9.992000000e-07 V_low
+ 9.992010000e-07 V_low
+ 9.993000000e-07 V_low
+ 9.993010000e-07 V_low
+ 9.994000000e-07 V_low
+ 9.994010000e-07 V_low
+ 9.995000000e-07 V_low
+ 9.995010000e-07 V_low
+ 9.996000000e-07 V_low
+ 9.996010000e-07 V_low
+ 9.997000000e-07 V_low
+ 9.997010000e-07 V_low
+ 9.998000000e-07 V_low
+ 9.998010000e-07 V_low
+ 9.999000000e-07 V_low
+ 9.999010000e-07 V_low
+ 1.000000000e-06 V_low
+ 1.000001000e-06 V_low
+ 1.000100000e-06 V_low
+ 1.000101000e-06 V_low
+ 1.000200000e-06 V_low
+ 1.000201000e-06 V_low
+ 1.000300000e-06 V_low
+ 1.000301000e-06 V_low
+ 1.000400000e-06 V_low
+ 1.000401000e-06 V_low
+ 1.000500000e-06 V_low
+ 1.000501000e-06 V_low
+ 1.000600000e-06 V_low
+ 1.000601000e-06 V_low
+ 1.000700000e-06 V_low
+ 1.000701000e-06 V_low
+ 1.000800000e-06 V_low
+ 1.000801000e-06 V_low
+ 1.000900000e-06 V_low
+ 
v2 b1 0 PWL
+ 1.000000000e-12 V_hig
+ 1.000000000e-09 V_hig
+ 1.001000000e-09 V_hig
+ 1.100000000e-09 V_hig
+ 1.101000000e-09 V_hig
+ 1.200000000e-09 V_hig
+ 1.201000000e-09 V_hig
+ 1.300000000e-09 V_hig
+ 1.301000000e-09 V_hig
+ 1.400000000e-09 V_hig
+ 1.401000000e-09 V_hig
+ 1.500000000e-09 V_hig
+ 1.501000000e-09 V_hig
+ 1.600000000e-09 V_hig
+ 1.601000000e-09 V_hig
+ 1.700000000e-09 V_hig
+ 1.701000000e-09 V_hig
+ 1.800000000e-09 V_hig
+ 1.801000000e-09 V_hig
+ 1.900000000e-09 V_hig
+ 1.901000000e-09 V_low
+ 2.000000000e-09 V_low
+ 2.001000000e-09 V_low
+ 2.100000000e-09 V_low
+ 2.101000000e-09 V_low
+ 2.200000000e-09 V_low
+ 2.201000000e-09 V_low
+ 2.300000000e-09 V_low
+ 2.301000000e-09 V_low
+ 2.400000000e-09 V_low
+ 2.401000000e-09 V_low
+ 2.500000000e-09 V_low
+ 2.501000000e-09 V_low
+ 2.600000000e-09 V_low
+ 2.601000000e-09 V_low
+ 2.700000000e-09 V_low
+ 2.701000000e-09 V_low
+ 2.800000000e-09 V_low
+ 2.801000000e-09 V_low
+ 2.900000000e-09 V_low
+ 2.901000000e-09 V_low
+ 3.000000000e-09 V_low
+ 3.001000000e-09 V_low
+ 3.100000000e-09 V_low
+ 3.101000000e-09 V_low
+ 3.200000000e-09 V_low
+ 3.201000000e-09 V_low
+ 3.300000000e-09 V_low
+ 3.301000000e-09 V_low
+ 3.400000000e-09 V_low
+ 3.401000000e-09 V_low
+ 3.500000000e-09 V_low
+ 3.501000000e-09 V_low
+ 3.600000000e-09 V_low
+ 3.601000000e-09 V_low
+ 3.700000000e-09 V_low
+ 3.701000000e-09 V_low
+ 3.800000000e-09 V_low
+ 3.801000000e-09 V_low
+ 3.900000000e-09 V_low
+ 3.901000000e-09 V_low
+ 4.000000000e-09 V_low
+ 4.001000000e-09 V_low
+ 4.100000000e-09 V_low
+ 4.101000000e-09 V_low
+ 4.200000000e-09 V_low
+ 4.201000000e-09 V_low
+ 4.300000000e-09 V_low
+ 4.301000000e-09 V_low
+ 4.400000000e-09 V_low
+ 4.401000000e-09 V_low
+ 4.500000000e-09 V_low
+ 4.501000000e-09 V_low
+ 4.600000000e-09 V_low
+ 4.601000000e-09 V_low
+ 4.700000000e-09 V_low
+ 4.701000000e-09 V_low
+ 4.800000000e-09 V_low
+ 4.801000000e-09 V_low
+ 4.900000000e-09 V_low
+ 4.901000000e-09 V_hig
+ 5.000000000e-09 V_hig
+ 5.001000000e-09 V_hig
+ 5.100000000e-09 V_hig
+ 5.101000000e-09 V_hig
+ 5.200000000e-09 V_hig
+ 5.201000000e-09 V_hig
+ 5.300000000e-09 V_hig
+ 5.301000000e-09 V_hig
+ 5.400000000e-09 V_hig
+ 5.401000000e-09 V_hig
+ 5.500000000e-09 V_hig
+ 5.501000000e-09 V_hig
+ 5.600000000e-09 V_hig
+ 5.601000000e-09 V_hig
+ 5.700000000e-09 V_hig
+ 5.701000000e-09 V_hig
+ 5.800000000e-09 V_hig
+ 5.801000000e-09 V_hig
+ 5.900000000e-09 V_hig
+ 5.901000000e-09 V_hig
+ 6.000000000e-09 V_hig
+ 6.001000000e-09 V_hig
+ 6.100000000e-09 V_hig
+ 6.101000000e-09 V_hig
+ 6.200000000e-09 V_hig
+ 6.201000000e-09 V_hig
+ 6.300000000e-09 V_hig
+ 6.301000000e-09 V_hig
+ 6.400000000e-09 V_hig
+ 6.401000000e-09 V_hig
+ 6.500000000e-09 V_hig
+ 6.501000000e-09 V_hig
+ 6.600000000e-09 V_hig
+ 6.601000000e-09 V_hig
+ 6.700000000e-09 V_hig
+ 6.701000000e-09 V_hig
+ 6.800000000e-09 V_hig
+ 6.801000000e-09 V_hig
+ 6.900000000e-09 V_hig
+ 6.901000000e-09 V_hig
+ 7.000000000e-09 V_hig
+ 7.001000000e-09 V_hig
+ 7.100000000e-09 V_hig
+ 7.101000000e-09 V_hig
+ 7.200000000e-09 V_hig
+ 7.201000000e-09 V_hig
+ 7.300000000e-09 V_hig
+ 7.301000000e-09 V_hig
+ 7.400000000e-09 V_hig
+ 7.401000000e-09 V_hig
+ 7.500000000e-09 V_hig
+ 7.501000000e-09 V_hig
+ 7.600000000e-09 V_hig
+ 7.601000000e-09 V_hig
+ 7.700000000e-09 V_hig
+ 7.701000000e-09 V_hig
+ 7.800000000e-09 V_hig
+ 7.801000000e-09 V_hig
+ 7.900000000e-09 V_hig
+ 7.901000000e-09 V_hig
+ 8.000000000e-09 V_hig
+ 8.001000000e-09 V_hig
+ 8.100000000e-09 V_hig
+ 8.101000000e-09 V_hig
+ 8.200000000e-09 V_hig
+ 8.201000000e-09 V_hig
+ 8.300000000e-09 V_hig
+ 8.301000000e-09 V_hig
+ 8.400000000e-09 V_hig
+ 8.401000000e-09 V_hig
+ 8.500000000e-09 V_hig
+ 8.501000000e-09 V_hig
+ 8.600000000e-09 V_hig
+ 8.601000000e-09 V_hig
+ 8.700000000e-09 V_hig
+ 8.701000000e-09 V_hig
+ 8.800000000e-09 V_hig
+ 8.801000000e-09 V_hig
+ 8.900000000e-09 V_hig
+ 8.901000000e-09 V_low
+ 9.000000000e-09 V_low
+ 9.001000000e-09 V_low
+ 9.100000000e-09 V_low
+ 9.101000000e-09 V_low
+ 9.200000000e-09 V_low
+ 9.201000000e-09 V_low
+ 9.300000000e-09 V_low
+ 9.301000000e-09 V_low
+ 9.400000000e-09 V_low
+ 9.401000000e-09 V_low
+ 9.500000000e-09 V_low
+ 9.501000000e-09 V_low
+ 9.600000000e-09 V_low
+ 9.601000000e-09 V_low
+ 9.700000000e-09 V_low
+ 9.701000000e-09 V_low
+ 9.800000000e-09 V_low
+ 9.801000000e-09 V_low
+ 9.900000000e-09 V_low
+ 9.901000000e-09 V_hig
+ 1.000000000e-08 V_hig
+ 1.000100000e-08 V_hig
+ 1.010000000e-08 V_hig
+ 1.010100000e-08 V_hig
+ 1.020000000e-08 V_hig
+ 1.020100000e-08 V_hig
+ 1.030000000e-08 V_hig
+ 1.030100000e-08 V_hig
+ 1.040000000e-08 V_hig
+ 1.040100000e-08 V_hig
+ 1.050000000e-08 V_hig
+ 1.050100000e-08 V_hig
+ 1.060000000e-08 V_hig
+ 1.060100000e-08 V_hig
+ 1.070000000e-08 V_hig
+ 1.070100000e-08 V_hig
+ 1.080000000e-08 V_hig
+ 1.080100000e-08 V_hig
+ 1.090000000e-08 V_hig
+ 1.090100000e-08 V_hig
+ 1.100000000e-08 V_hig
+ 1.100100000e-08 V_hig
+ 1.110000000e-08 V_hig
+ 1.110100000e-08 V_hig
+ 1.120000000e-08 V_hig
+ 1.120100000e-08 V_hig
+ 1.130000000e-08 V_hig
+ 1.130100000e-08 V_hig
+ 1.140000000e-08 V_hig
+ 1.140100000e-08 V_hig
+ 1.150000000e-08 V_hig
+ 1.150100000e-08 V_hig
+ 1.160000000e-08 V_hig
+ 1.160100000e-08 V_hig
+ 1.170000000e-08 V_hig
+ 1.170100000e-08 V_hig
+ 1.180000000e-08 V_hig
+ 1.180100000e-08 V_hig
+ 1.190000000e-08 V_hig
+ 1.190100000e-08 V_hig
+ 1.200000000e-08 V_hig
+ 1.200100000e-08 V_hig
+ 1.210000000e-08 V_hig
+ 1.210100000e-08 V_hig
+ 1.220000000e-08 V_hig
+ 1.220100000e-08 V_hig
+ 1.230000000e-08 V_hig
+ 1.230100000e-08 V_hig
+ 1.240000000e-08 V_hig
+ 1.240100000e-08 V_hig
+ 1.250000000e-08 V_hig
+ 1.250100000e-08 V_hig
+ 1.260000000e-08 V_hig
+ 1.260100000e-08 V_hig
+ 1.270000000e-08 V_hig
+ 1.270100000e-08 V_hig
+ 1.280000000e-08 V_hig
+ 1.280100000e-08 V_hig
+ 1.290000000e-08 V_hig
+ 1.290100000e-08 V_hig
+ 1.300000000e-08 V_hig
+ 1.300100000e-08 V_hig
+ 1.310000000e-08 V_hig
+ 1.310100000e-08 V_hig
+ 1.320000000e-08 V_hig
+ 1.320100000e-08 V_hig
+ 1.330000000e-08 V_hig
+ 1.330100000e-08 V_hig
+ 1.340000000e-08 V_hig
+ 1.340100000e-08 V_hig
+ 1.350000000e-08 V_hig
+ 1.350100000e-08 V_hig
+ 1.360000000e-08 V_hig
+ 1.360100000e-08 V_hig
+ 1.370000000e-08 V_hig
+ 1.370100000e-08 V_hig
+ 1.380000000e-08 V_hig
+ 1.380100000e-08 V_hig
+ 1.390000000e-08 V_hig
+ 1.390100000e-08 V_low
+ 1.400000000e-08 V_low
+ 1.400100000e-08 V_low
+ 1.410000000e-08 V_low
+ 1.410100000e-08 V_low
+ 1.420000000e-08 V_low
+ 1.420100000e-08 V_low
+ 1.430000000e-08 V_low
+ 1.430100000e-08 V_low
+ 1.440000000e-08 V_low
+ 1.440100000e-08 V_low
+ 1.450000000e-08 V_low
+ 1.450100000e-08 V_low
+ 1.460000000e-08 V_low
+ 1.460100000e-08 V_low
+ 1.470000000e-08 V_low
+ 1.470100000e-08 V_low
+ 1.480000000e-08 V_low
+ 1.480100000e-08 V_low
+ 1.490000000e-08 V_low
+ 1.490100000e-08 V_hig
+ 1.500000000e-08 V_hig
+ 1.500100000e-08 V_hig
+ 1.510000000e-08 V_hig
+ 1.510100000e-08 V_hig
+ 1.520000000e-08 V_hig
+ 1.520100000e-08 V_hig
+ 1.530000000e-08 V_hig
+ 1.530100000e-08 V_hig
+ 1.540000000e-08 V_hig
+ 1.540100000e-08 V_hig
+ 1.550000000e-08 V_hig
+ 1.550100000e-08 V_hig
+ 1.560000000e-08 V_hig
+ 1.560100000e-08 V_hig
+ 1.570000000e-08 V_hig
+ 1.570100000e-08 V_hig
+ 1.580000000e-08 V_hig
+ 1.580100000e-08 V_hig
+ 1.590000000e-08 V_hig
+ 1.590100000e-08 V_low
+ 1.600000000e-08 V_low
+ 1.600100000e-08 V_low
+ 1.610000000e-08 V_low
+ 1.610100000e-08 V_low
+ 1.620000000e-08 V_low
+ 1.620100000e-08 V_low
+ 1.630000000e-08 V_low
+ 1.630100000e-08 V_low
+ 1.640000000e-08 V_low
+ 1.640100000e-08 V_low
+ 1.650000000e-08 V_low
+ 1.650100000e-08 V_low
+ 1.660000000e-08 V_low
+ 1.660100000e-08 V_low
+ 1.670000000e-08 V_low
+ 1.670100000e-08 V_low
+ 1.680000000e-08 V_low
+ 1.680100000e-08 V_low
+ 1.690000000e-08 V_low
+ 1.690100000e-08 V_low
+ 1.700000000e-08 V_low
+ 1.700100000e-08 V_low
+ 1.710000000e-08 V_low
+ 1.710100000e-08 V_low
+ 1.720000000e-08 V_low
+ 1.720100000e-08 V_low
+ 1.730000000e-08 V_low
+ 1.730100000e-08 V_low
+ 1.740000000e-08 V_low
+ 1.740100000e-08 V_low
+ 1.750000000e-08 V_low
+ 1.750100000e-08 V_low
+ 1.760000000e-08 V_low
+ 1.760100000e-08 V_low
+ 1.770000000e-08 V_low
+ 1.770100000e-08 V_low
+ 1.780000000e-08 V_low
+ 1.780100000e-08 V_low
+ 1.790000000e-08 V_low
+ 1.790100000e-08 V_hig
+ 1.800000000e-08 V_hig
+ 1.800100000e-08 V_hig
+ 1.810000000e-08 V_hig
+ 1.810100000e-08 V_hig
+ 1.820000000e-08 V_hig
+ 1.820100000e-08 V_hig
+ 1.830000000e-08 V_hig
+ 1.830100000e-08 V_hig
+ 1.840000000e-08 V_hig
+ 1.840100000e-08 V_hig
+ 1.850000000e-08 V_hig
+ 1.850100000e-08 V_hig
+ 1.860000000e-08 V_hig
+ 1.860100000e-08 V_hig
+ 1.870000000e-08 V_hig
+ 1.870100000e-08 V_hig
+ 1.880000000e-08 V_hig
+ 1.880100000e-08 V_hig
+ 1.890000000e-08 V_hig
+ 1.890100000e-08 V_low
+ 1.900000000e-08 V_low
+ 1.900100000e-08 V_low
+ 1.910000000e-08 V_low
+ 1.910100000e-08 V_low
+ 1.920000000e-08 V_low
+ 1.920100000e-08 V_low
+ 1.930000000e-08 V_low
+ 1.930100000e-08 V_low
+ 1.940000000e-08 V_low
+ 1.940100000e-08 V_low
+ 1.950000000e-08 V_low
+ 1.950100000e-08 V_low
+ 1.960000000e-08 V_low
+ 1.960100000e-08 V_low
+ 1.970000000e-08 V_low
+ 1.970100000e-08 V_low
+ 1.980000000e-08 V_low
+ 1.980100000e-08 V_low
+ 1.990000000e-08 V_low
+ 1.990100000e-08 V_low
+ 2.000000000e-08 V_low
+ 2.000100000e-08 V_low
+ 2.010000000e-08 V_low
+ 2.010100000e-08 V_low
+ 2.020000000e-08 V_low
+ 2.020100000e-08 V_low
+ 2.030000000e-08 V_low
+ 2.030100000e-08 V_low
+ 2.040000000e-08 V_low
+ 2.040100000e-08 V_low
+ 2.050000000e-08 V_low
+ 2.050100000e-08 V_low
+ 2.060000000e-08 V_low
+ 2.060100000e-08 V_low
+ 2.070000000e-08 V_low
+ 2.070100000e-08 V_low
+ 2.080000000e-08 V_low
+ 2.080100000e-08 V_low
+ 2.090000000e-08 V_low
+ 2.090100000e-08 V_low
+ 2.100000000e-08 V_low
+ 2.100100000e-08 V_low
+ 2.110000000e-08 V_low
+ 2.110100000e-08 V_low
+ 2.120000000e-08 V_low
+ 2.120100000e-08 V_low
+ 2.130000000e-08 V_low
+ 2.130100000e-08 V_low
+ 2.140000000e-08 V_low
+ 2.140100000e-08 V_low
+ 2.150000000e-08 V_low
+ 2.150100000e-08 V_low
+ 2.160000000e-08 V_low
+ 2.160100000e-08 V_low
+ 2.170000000e-08 V_low
+ 2.170100000e-08 V_low
+ 2.180000000e-08 V_low
+ 2.180100000e-08 V_low
+ 2.190000000e-08 V_low
+ 2.190100000e-08 V_low
+ 2.200000000e-08 V_low
+ 2.200100000e-08 V_low
+ 2.210000000e-08 V_low
+ 2.210100000e-08 V_low
+ 2.220000000e-08 V_low
+ 2.220100000e-08 V_low
+ 2.230000000e-08 V_low
+ 2.230100000e-08 V_low
+ 2.240000000e-08 V_low
+ 2.240100000e-08 V_low
+ 2.250000000e-08 V_low
+ 2.250100000e-08 V_low
+ 2.260000000e-08 V_low
+ 2.260100000e-08 V_low
+ 2.270000000e-08 V_low
+ 2.270100000e-08 V_low
+ 2.280000000e-08 V_low
+ 2.280100000e-08 V_low
+ 2.290000000e-08 V_low
+ 2.290100000e-08 V_low
+ 2.300000000e-08 V_low
+ 2.300100000e-08 V_low
+ 2.310000000e-08 V_low
+ 2.310100000e-08 V_low
+ 2.320000000e-08 V_low
+ 2.320100000e-08 V_low
+ 2.330000000e-08 V_low
+ 2.330100000e-08 V_low
+ 2.340000000e-08 V_low
+ 2.340100000e-08 V_low
+ 2.350000000e-08 V_low
+ 2.350100000e-08 V_low
+ 2.360000000e-08 V_low
+ 2.360100000e-08 V_low
+ 2.370000000e-08 V_low
+ 2.370100000e-08 V_low
+ 2.380000000e-08 V_low
+ 2.380100000e-08 V_low
+ 2.390000000e-08 V_low
+ 2.390100000e-08 V_hig
+ 2.400000000e-08 V_hig
+ 2.400100000e-08 V_hig
+ 2.410000000e-08 V_hig
+ 2.410100000e-08 V_hig
+ 2.420000000e-08 V_hig
+ 2.420100000e-08 V_hig
+ 2.430000000e-08 V_hig
+ 2.430100000e-08 V_hig
+ 2.440000000e-08 V_hig
+ 2.440100000e-08 V_hig
+ 2.450000000e-08 V_hig
+ 2.450100000e-08 V_hig
+ 2.460000000e-08 V_hig
+ 2.460100000e-08 V_hig
+ 2.470000000e-08 V_hig
+ 2.470100000e-08 V_hig
+ 2.480000000e-08 V_hig
+ 2.480100000e-08 V_hig
+ 2.490000000e-08 V_hig
+ 2.490100000e-08 V_hig
+ 2.500000000e-08 V_hig
+ 2.500100000e-08 V_hig
+ 2.510000000e-08 V_hig
+ 2.510100000e-08 V_hig
+ 2.520000000e-08 V_hig
+ 2.520100000e-08 V_hig
+ 2.530000000e-08 V_hig
+ 2.530100000e-08 V_hig
+ 2.540000000e-08 V_hig
+ 2.540100000e-08 V_hig
+ 2.550000000e-08 V_hig
+ 2.550100000e-08 V_hig
+ 2.560000000e-08 V_hig
+ 2.560100000e-08 V_hig
+ 2.570000000e-08 V_hig
+ 2.570100000e-08 V_hig
+ 2.580000000e-08 V_hig
+ 2.580100000e-08 V_hig
+ 2.590000000e-08 V_hig
+ 2.590100000e-08 V_hig
+ 2.600000000e-08 V_hig
+ 2.600100000e-08 V_hig
+ 2.610000000e-08 V_hig
+ 2.610100000e-08 V_hig
+ 2.620000000e-08 V_hig
+ 2.620100000e-08 V_hig
+ 2.630000000e-08 V_hig
+ 2.630100000e-08 V_hig
+ 2.640000000e-08 V_hig
+ 2.640100000e-08 V_hig
+ 2.650000000e-08 V_hig
+ 2.650100000e-08 V_hig
+ 2.660000000e-08 V_hig
+ 2.660100000e-08 V_hig
+ 2.670000000e-08 V_hig
+ 2.670100000e-08 V_hig
+ 2.680000000e-08 V_hig
+ 2.680100000e-08 V_hig
+ 2.690000000e-08 V_hig
+ 2.690100000e-08 V_low
+ 2.700000000e-08 V_low
+ 2.700100000e-08 V_low
+ 2.710000000e-08 V_low
+ 2.710100000e-08 V_low
+ 2.720000000e-08 V_low
+ 2.720100000e-08 V_low
+ 2.730000000e-08 V_low
+ 2.730100000e-08 V_low
+ 2.740000000e-08 V_low
+ 2.740100000e-08 V_low
+ 2.750000000e-08 V_low
+ 2.750100000e-08 V_low
+ 2.760000000e-08 V_low
+ 2.760100000e-08 V_low
+ 2.770000000e-08 V_low
+ 2.770100000e-08 V_low
+ 2.780000000e-08 V_low
+ 2.780100000e-08 V_low
+ 2.790000000e-08 V_low
+ 2.790100000e-08 V_hig
+ 2.800000000e-08 V_hig
+ 2.800100000e-08 V_hig
+ 2.810000000e-08 V_hig
+ 2.810100000e-08 V_hig
+ 2.820000000e-08 V_hig
+ 2.820100000e-08 V_hig
+ 2.830000000e-08 V_hig
+ 2.830100000e-08 V_hig
+ 2.840000000e-08 V_hig
+ 2.840100000e-08 V_hig
+ 2.850000000e-08 V_hig
+ 2.850100000e-08 V_hig
+ 2.860000000e-08 V_hig
+ 2.860100000e-08 V_hig
+ 2.870000000e-08 V_hig
+ 2.870100000e-08 V_hig
+ 2.880000000e-08 V_hig
+ 2.880100000e-08 V_hig
+ 2.890000000e-08 V_hig
+ 2.890100000e-08 V_low
+ 2.900000000e-08 V_low
+ 2.900100000e-08 V_low
+ 2.910000000e-08 V_low
+ 2.910100000e-08 V_low
+ 2.920000000e-08 V_low
+ 2.920100000e-08 V_low
+ 2.930000000e-08 V_low
+ 2.930100000e-08 V_low
+ 2.940000000e-08 V_low
+ 2.940100000e-08 V_low
+ 2.950000000e-08 V_low
+ 2.950100000e-08 V_low
+ 2.960000000e-08 V_low
+ 2.960100000e-08 V_low
+ 2.970000000e-08 V_low
+ 2.970100000e-08 V_low
+ 2.980000000e-08 V_low
+ 2.980100000e-08 V_low
+ 2.990000000e-08 V_low
+ 2.990100000e-08 V_hig
+ 3.000000000e-08 V_hig
+ 3.000100000e-08 V_hig
+ 3.010000000e-08 V_hig
+ 3.010100000e-08 V_hig
+ 3.020000000e-08 V_hig
+ 3.020100000e-08 V_hig
+ 3.030000000e-08 V_hig
+ 3.030100000e-08 V_hig
+ 3.040000000e-08 V_hig
+ 3.040100000e-08 V_hig
+ 3.050000000e-08 V_hig
+ 3.050100000e-08 V_hig
+ 3.060000000e-08 V_hig
+ 3.060100000e-08 V_hig
+ 3.070000000e-08 V_hig
+ 3.070100000e-08 V_hig
+ 3.080000000e-08 V_hig
+ 3.080100000e-08 V_hig
+ 3.090000000e-08 V_hig
+ 3.090100000e-08 V_hig
+ 3.100000000e-08 V_hig
+ 3.100100000e-08 V_hig
+ 3.110000000e-08 V_hig
+ 3.110100000e-08 V_hig
+ 3.120000000e-08 V_hig
+ 3.120100000e-08 V_hig
+ 3.130000000e-08 V_hig
+ 3.130100000e-08 V_hig
+ 3.140000000e-08 V_hig
+ 3.140100000e-08 V_hig
+ 3.150000000e-08 V_hig
+ 3.150100000e-08 V_hig
+ 3.160000000e-08 V_hig
+ 3.160100000e-08 V_hig
+ 3.170000000e-08 V_hig
+ 3.170100000e-08 V_hig
+ 3.180000000e-08 V_hig
+ 3.180100000e-08 V_hig
+ 3.190000000e-08 V_hig
+ 3.190100000e-08 V_low
+ 3.200000000e-08 V_low
+ 3.200100000e-08 V_low
+ 3.210000000e-08 V_low
+ 3.210100000e-08 V_low
+ 3.220000000e-08 V_low
+ 3.220100000e-08 V_low
+ 3.230000000e-08 V_low
+ 3.230100000e-08 V_low
+ 3.240000000e-08 V_low
+ 3.240100000e-08 V_low
+ 3.250000000e-08 V_low
+ 3.250100000e-08 V_low
+ 3.260000000e-08 V_low
+ 3.260100000e-08 V_low
+ 3.270000000e-08 V_low
+ 3.270100000e-08 V_low
+ 3.280000000e-08 V_low
+ 3.280100000e-08 V_low
+ 3.290000000e-08 V_low
+ 3.290100000e-08 V_hig
+ 3.300000000e-08 V_hig
+ 3.300100000e-08 V_hig
+ 3.310000000e-08 V_hig
+ 3.310100000e-08 V_hig
+ 3.320000000e-08 V_hig
+ 3.320100000e-08 V_hig
+ 3.330000000e-08 V_hig
+ 3.330100000e-08 V_hig
+ 3.340000000e-08 V_hig
+ 3.340100000e-08 V_hig
+ 3.350000000e-08 V_hig
+ 3.350100000e-08 V_hig
+ 3.360000000e-08 V_hig
+ 3.360100000e-08 V_hig
+ 3.370000000e-08 V_hig
+ 3.370100000e-08 V_hig
+ 3.380000000e-08 V_hig
+ 3.380100000e-08 V_hig
+ 3.390000000e-08 V_hig
+ 3.390100000e-08 V_low
+ 3.400000000e-08 V_low
+ 3.400100000e-08 V_low
+ 3.410000000e-08 V_low
+ 3.410100000e-08 V_low
+ 3.420000000e-08 V_low
+ 3.420100000e-08 V_low
+ 3.430000000e-08 V_low
+ 3.430100000e-08 V_low
+ 3.440000000e-08 V_low
+ 3.440100000e-08 V_low
+ 3.450000000e-08 V_low
+ 3.450100000e-08 V_low
+ 3.460000000e-08 V_low
+ 3.460100000e-08 V_low
+ 3.470000000e-08 V_low
+ 3.470100000e-08 V_low
+ 3.480000000e-08 V_low
+ 3.480100000e-08 V_low
+ 3.490000000e-08 V_low
+ 3.490100000e-08 V_low
+ 3.500000000e-08 V_low
+ 3.500100000e-08 V_low
+ 3.510000000e-08 V_low
+ 3.510100000e-08 V_low
+ 3.520000000e-08 V_low
+ 3.520100000e-08 V_low
+ 3.530000000e-08 V_low
+ 3.530100000e-08 V_low
+ 3.540000000e-08 V_low
+ 3.540100000e-08 V_low
+ 3.550000000e-08 V_low
+ 3.550100000e-08 V_low
+ 3.560000000e-08 V_low
+ 3.560100000e-08 V_low
+ 3.570000000e-08 V_low
+ 3.570100000e-08 V_low
+ 3.580000000e-08 V_low
+ 3.580100000e-08 V_low
+ 3.590000000e-08 V_low
+ 3.590100000e-08 V_hig
+ 3.600000000e-08 V_hig
+ 3.600100000e-08 V_hig
+ 3.610000000e-08 V_hig
+ 3.610100000e-08 V_hig
+ 3.620000000e-08 V_hig
+ 3.620100000e-08 V_hig
+ 3.630000000e-08 V_hig
+ 3.630100000e-08 V_hig
+ 3.640000000e-08 V_hig
+ 3.640100000e-08 V_hig
+ 3.650000000e-08 V_hig
+ 3.650100000e-08 V_hig
+ 3.660000000e-08 V_hig
+ 3.660100000e-08 V_hig
+ 3.670000000e-08 V_hig
+ 3.670100000e-08 V_hig
+ 3.680000000e-08 V_hig
+ 3.680100000e-08 V_hig
+ 3.690000000e-08 V_hig
+ 3.690100000e-08 V_hig
+ 3.700000000e-08 V_hig
+ 3.700100000e-08 V_hig
+ 3.710000000e-08 V_hig
+ 3.710100000e-08 V_hig
+ 3.720000000e-08 V_hig
+ 3.720100000e-08 V_hig
+ 3.730000000e-08 V_hig
+ 3.730100000e-08 V_hig
+ 3.740000000e-08 V_hig
+ 3.740100000e-08 V_hig
+ 3.750000000e-08 V_hig
+ 3.750100000e-08 V_hig
+ 3.760000000e-08 V_hig
+ 3.760100000e-08 V_hig
+ 3.770000000e-08 V_hig
+ 3.770100000e-08 V_hig
+ 3.780000000e-08 V_hig
+ 3.780100000e-08 V_hig
+ 3.790000000e-08 V_hig
+ 3.790100000e-08 V_low
+ 3.800000000e-08 V_low
+ 3.800100000e-08 V_low
+ 3.810000000e-08 V_low
+ 3.810100000e-08 V_low
+ 3.820000000e-08 V_low
+ 3.820100000e-08 V_low
+ 3.830000000e-08 V_low
+ 3.830100000e-08 V_low
+ 3.840000000e-08 V_low
+ 3.840100000e-08 V_low
+ 3.850000000e-08 V_low
+ 3.850100000e-08 V_low
+ 3.860000000e-08 V_low
+ 3.860100000e-08 V_low
+ 3.870000000e-08 V_low
+ 3.870100000e-08 V_low
+ 3.880000000e-08 V_low
+ 3.880100000e-08 V_low
+ 3.890000000e-08 V_low
+ 3.890100000e-08 V_hig
+ 3.900000000e-08 V_hig
+ 3.900100000e-08 V_hig
+ 3.910000000e-08 V_hig
+ 3.910100000e-08 V_hig
+ 3.920000000e-08 V_hig
+ 3.920100000e-08 V_hig
+ 3.930000000e-08 V_hig
+ 3.930100000e-08 V_hig
+ 3.940000000e-08 V_hig
+ 3.940100000e-08 V_hig
+ 3.950000000e-08 V_hig
+ 3.950100000e-08 V_hig
+ 3.960000000e-08 V_hig
+ 3.960100000e-08 V_hig
+ 3.970000000e-08 V_hig
+ 3.970100000e-08 V_hig
+ 3.980000000e-08 V_hig
+ 3.980100000e-08 V_hig
+ 3.990000000e-08 V_hig
+ 3.990100000e-08 V_hig
+ 4.000000000e-08 V_hig
+ 4.000100000e-08 V_hig
+ 4.010000000e-08 V_hig
+ 4.010100000e-08 V_hig
+ 4.020000000e-08 V_hig
+ 4.020100000e-08 V_hig
+ 4.030000000e-08 V_hig
+ 4.030100000e-08 V_hig
+ 4.040000000e-08 V_hig
+ 4.040100000e-08 V_hig
+ 4.050000000e-08 V_hig
+ 4.050100000e-08 V_hig
+ 4.060000000e-08 V_hig
+ 4.060100000e-08 V_hig
+ 4.070000000e-08 V_hig
+ 4.070100000e-08 V_hig
+ 4.080000000e-08 V_hig
+ 4.080100000e-08 V_hig
+ 4.090000000e-08 V_hig
+ 4.090100000e-08 V_hig
+ 4.100000000e-08 V_hig
+ 4.100100000e-08 V_hig
+ 4.110000000e-08 V_hig
+ 4.110100000e-08 V_hig
+ 4.120000000e-08 V_hig
+ 4.120100000e-08 V_hig
+ 4.130000000e-08 V_hig
+ 4.130100000e-08 V_hig
+ 4.140000000e-08 V_hig
+ 4.140100000e-08 V_hig
+ 4.150000000e-08 V_hig
+ 4.150100000e-08 V_hig
+ 4.160000000e-08 V_hig
+ 4.160100000e-08 V_hig
+ 4.170000000e-08 V_hig
+ 4.170100000e-08 V_hig
+ 4.180000000e-08 V_hig
+ 4.180100000e-08 V_hig
+ 4.190000000e-08 V_hig
+ 4.190100000e-08 V_hig
+ 4.200000000e-08 V_hig
+ 4.200100000e-08 V_hig
+ 4.210000000e-08 V_hig
+ 4.210100000e-08 V_hig
+ 4.220000000e-08 V_hig
+ 4.220100000e-08 V_hig
+ 4.230000000e-08 V_hig
+ 4.230100000e-08 V_hig
+ 4.240000000e-08 V_hig
+ 4.240100000e-08 V_hig
+ 4.250000000e-08 V_hig
+ 4.250100000e-08 V_hig
+ 4.260000000e-08 V_hig
+ 4.260100000e-08 V_hig
+ 4.270000000e-08 V_hig
+ 4.270100000e-08 V_hig
+ 4.280000000e-08 V_hig
+ 4.280100000e-08 V_hig
+ 4.290000000e-08 V_hig
+ 4.290100000e-08 V_low
+ 4.300000000e-08 V_low
+ 4.300100000e-08 V_low
+ 4.310000000e-08 V_low
+ 4.310100000e-08 V_low
+ 4.320000000e-08 V_low
+ 4.320100000e-08 V_low
+ 4.330000000e-08 V_low
+ 4.330100000e-08 V_low
+ 4.340000000e-08 V_low
+ 4.340100000e-08 V_low
+ 4.350000000e-08 V_low
+ 4.350100000e-08 V_low
+ 4.360000000e-08 V_low
+ 4.360100000e-08 V_low
+ 4.370000000e-08 V_low
+ 4.370100000e-08 V_low
+ 4.380000000e-08 V_low
+ 4.380100000e-08 V_low
+ 4.390000000e-08 V_low
+ 4.390100000e-08 V_low
+ 4.400000000e-08 V_low
+ 4.400100000e-08 V_low
+ 4.410000000e-08 V_low
+ 4.410100000e-08 V_low
+ 4.420000000e-08 V_low
+ 4.420100000e-08 V_low
+ 4.430000000e-08 V_low
+ 4.430100000e-08 V_low
+ 4.440000000e-08 V_low
+ 4.440100000e-08 V_low
+ 4.450000000e-08 V_low
+ 4.450100000e-08 V_low
+ 4.460000000e-08 V_low
+ 4.460100000e-08 V_low
+ 4.470000000e-08 V_low
+ 4.470100000e-08 V_low
+ 4.480000000e-08 V_low
+ 4.480100000e-08 V_low
+ 4.490000000e-08 V_low
+ 4.490100000e-08 V_hig
+ 4.500000000e-08 V_hig
+ 4.500100000e-08 V_hig
+ 4.510000000e-08 V_hig
+ 4.510100000e-08 V_hig
+ 4.520000000e-08 V_hig
+ 4.520100000e-08 V_hig
+ 4.530000000e-08 V_hig
+ 4.530100000e-08 V_hig
+ 4.540000000e-08 V_hig
+ 4.540100000e-08 V_hig
+ 4.550000000e-08 V_hig
+ 4.550100000e-08 V_hig
+ 4.560000000e-08 V_hig
+ 4.560100000e-08 V_hig
+ 4.570000000e-08 V_hig
+ 4.570100000e-08 V_hig
+ 4.580000000e-08 V_hig
+ 4.580100000e-08 V_hig
+ 4.590000000e-08 V_hig
+ 4.590100000e-08 V_hig
+ 4.600000000e-08 V_hig
+ 4.600100000e-08 V_hig
+ 4.610000000e-08 V_hig
+ 4.610100000e-08 V_hig
+ 4.620000000e-08 V_hig
+ 4.620100000e-08 V_hig
+ 4.630000000e-08 V_hig
+ 4.630100000e-08 V_hig
+ 4.640000000e-08 V_hig
+ 4.640100000e-08 V_hig
+ 4.650000000e-08 V_hig
+ 4.650100000e-08 V_hig
+ 4.660000000e-08 V_hig
+ 4.660100000e-08 V_hig
+ 4.670000000e-08 V_hig
+ 4.670100000e-08 V_hig
+ 4.680000000e-08 V_hig
+ 4.680100000e-08 V_hig
+ 4.690000000e-08 V_hig
+ 4.690100000e-08 V_low
+ 4.700000000e-08 V_low
+ 4.700100000e-08 V_low
+ 4.710000000e-08 V_low
+ 4.710100000e-08 V_low
+ 4.720000000e-08 V_low
+ 4.720100000e-08 V_low
+ 4.730000000e-08 V_low
+ 4.730100000e-08 V_low
+ 4.740000000e-08 V_low
+ 4.740100000e-08 V_low
+ 4.750000000e-08 V_low
+ 4.750100000e-08 V_low
+ 4.760000000e-08 V_low
+ 4.760100000e-08 V_low
+ 4.770000000e-08 V_low
+ 4.770100000e-08 V_low
+ 4.780000000e-08 V_low
+ 4.780100000e-08 V_low
+ 4.790000000e-08 V_low
+ 4.790100000e-08 V_low
+ 4.800000000e-08 V_low
+ 4.800100000e-08 V_low
+ 4.810000000e-08 V_low
+ 4.810100000e-08 V_low
+ 4.820000000e-08 V_low
+ 4.820100000e-08 V_low
+ 4.830000000e-08 V_low
+ 4.830100000e-08 V_low
+ 4.840000000e-08 V_low
+ 4.840100000e-08 V_low
+ 4.850000000e-08 V_low
+ 4.850100000e-08 V_low
+ 4.860000000e-08 V_low
+ 4.860100000e-08 V_low
+ 4.870000000e-08 V_low
+ 4.870100000e-08 V_low
+ 4.880000000e-08 V_low
+ 4.880100000e-08 V_low
+ 4.890000000e-08 V_low
+ 4.890100000e-08 V_low
+ 4.900000000e-08 V_low
+ 4.900100000e-08 V_low
+ 4.910000000e-08 V_low
+ 4.910100000e-08 V_low
+ 4.920000000e-08 V_low
+ 4.920100000e-08 V_low
+ 4.930000000e-08 V_low
+ 4.930100000e-08 V_low
+ 4.940000000e-08 V_low
+ 4.940100000e-08 V_low
+ 4.950000000e-08 V_low
+ 4.950100000e-08 V_low
+ 4.960000000e-08 V_low
+ 4.960100000e-08 V_low
+ 4.970000000e-08 V_low
+ 4.970100000e-08 V_low
+ 4.980000000e-08 V_low
+ 4.980100000e-08 V_low
+ 4.990000000e-08 V_low
+ 4.990100000e-08 V_low
+ 5.000000000e-08 V_low
+ 5.000100000e-08 V_low
+ 5.010000000e-08 V_low
+ 5.010100000e-08 V_low
+ 5.020000000e-08 V_low
+ 5.020100000e-08 V_low
+ 5.030000000e-08 V_low
+ 5.030100000e-08 V_low
+ 5.040000000e-08 V_low
+ 5.040100000e-08 V_low
+ 5.050000000e-08 V_low
+ 5.050100000e-08 V_low
+ 5.060000000e-08 V_low
+ 5.060100000e-08 V_low
+ 5.070000000e-08 V_low
+ 5.070100000e-08 V_low
+ 5.080000000e-08 V_low
+ 5.080100000e-08 V_low
+ 5.090000000e-08 V_low
+ 5.090100000e-08 V_low
+ 5.100000000e-08 V_low
+ 5.100100000e-08 V_low
+ 5.110000000e-08 V_low
+ 5.110100000e-08 V_low
+ 5.120000000e-08 V_low
+ 5.120100000e-08 V_low
+ 5.130000000e-08 V_low
+ 5.130100000e-08 V_low
+ 5.140000000e-08 V_low
+ 5.140100000e-08 V_low
+ 5.150000000e-08 V_low
+ 5.150100000e-08 V_low
+ 5.160000000e-08 V_low
+ 5.160100000e-08 V_low
+ 5.170000000e-08 V_low
+ 5.170100000e-08 V_low
+ 5.180000000e-08 V_low
+ 5.180100000e-08 V_low
+ 5.190000000e-08 V_low
+ 5.190100000e-08 V_low
+ 5.200000000e-08 V_low
+ 5.200100000e-08 V_low
+ 5.210000000e-08 V_low
+ 5.210100000e-08 V_low
+ 5.220000000e-08 V_low
+ 5.220100000e-08 V_low
+ 5.230000000e-08 V_low
+ 5.230100000e-08 V_low
+ 5.240000000e-08 V_low
+ 5.240100000e-08 V_low
+ 5.250000000e-08 V_low
+ 5.250100000e-08 V_low
+ 5.260000000e-08 V_low
+ 5.260100000e-08 V_low
+ 5.270000000e-08 V_low
+ 5.270100000e-08 V_low
+ 5.280000000e-08 V_low
+ 5.280100000e-08 V_low
+ 5.290000000e-08 V_low
+ 5.290100000e-08 V_low
+ 5.300000000e-08 V_low
+ 5.300100000e-08 V_low
+ 5.310000000e-08 V_low
+ 5.310100000e-08 V_low
+ 5.320000000e-08 V_low
+ 5.320100000e-08 V_low
+ 5.330000000e-08 V_low
+ 5.330100000e-08 V_low
+ 5.340000000e-08 V_low
+ 5.340100000e-08 V_low
+ 5.350000000e-08 V_low
+ 5.350100000e-08 V_low
+ 5.360000000e-08 V_low
+ 5.360100000e-08 V_low
+ 5.370000000e-08 V_low
+ 5.370100000e-08 V_low
+ 5.380000000e-08 V_low
+ 5.380100000e-08 V_low
+ 5.390000000e-08 V_low
+ 5.390100000e-08 V_hig
+ 5.400000000e-08 V_hig
+ 5.400100000e-08 V_hig
+ 5.410000000e-08 V_hig
+ 5.410100000e-08 V_hig
+ 5.420000000e-08 V_hig
+ 5.420100000e-08 V_hig
+ 5.430000000e-08 V_hig
+ 5.430100000e-08 V_hig
+ 5.440000000e-08 V_hig
+ 5.440100000e-08 V_hig
+ 5.450000000e-08 V_hig
+ 5.450100000e-08 V_hig
+ 5.460000000e-08 V_hig
+ 5.460100000e-08 V_hig
+ 5.470000000e-08 V_hig
+ 5.470100000e-08 V_hig
+ 5.480000000e-08 V_hig
+ 5.480100000e-08 V_hig
+ 5.490000000e-08 V_hig
+ 5.490100000e-08 V_low
+ 5.500000000e-08 V_low
+ 5.500100000e-08 V_low
+ 5.510000000e-08 V_low
+ 5.510100000e-08 V_low
+ 5.520000000e-08 V_low
+ 5.520100000e-08 V_low
+ 5.530000000e-08 V_low
+ 5.530100000e-08 V_low
+ 5.540000000e-08 V_low
+ 5.540100000e-08 V_low
+ 5.550000000e-08 V_low
+ 5.550100000e-08 V_low
+ 5.560000000e-08 V_low
+ 5.560100000e-08 V_low
+ 5.570000000e-08 V_low
+ 5.570100000e-08 V_low
+ 5.580000000e-08 V_low
+ 5.580100000e-08 V_low
+ 5.590000000e-08 V_low
+ 5.590100000e-08 V_low
+ 5.600000000e-08 V_low
+ 5.600100000e-08 V_low
+ 5.610000000e-08 V_low
+ 5.610100000e-08 V_low
+ 5.620000000e-08 V_low
+ 5.620100000e-08 V_low
+ 5.630000000e-08 V_low
+ 5.630100000e-08 V_low
+ 5.640000000e-08 V_low
+ 5.640100000e-08 V_low
+ 5.650000000e-08 V_low
+ 5.650100000e-08 V_low
+ 5.660000000e-08 V_low
+ 5.660100000e-08 V_low
+ 5.670000000e-08 V_low
+ 5.670100000e-08 V_low
+ 5.680000000e-08 V_low
+ 5.680100000e-08 V_low
+ 5.690000000e-08 V_low
+ 5.690100000e-08 V_low
+ 5.700000000e-08 V_low
+ 5.700100000e-08 V_low
+ 5.710000000e-08 V_low
+ 5.710100000e-08 V_low
+ 5.720000000e-08 V_low
+ 5.720100000e-08 V_low
+ 5.730000000e-08 V_low
+ 5.730100000e-08 V_low
+ 5.740000000e-08 V_low
+ 5.740100000e-08 V_low
+ 5.750000000e-08 V_low
+ 5.750100000e-08 V_low
+ 5.760000000e-08 V_low
+ 5.760100000e-08 V_low
+ 5.770000000e-08 V_low
+ 5.770100000e-08 V_low
+ 5.780000000e-08 V_low
+ 5.780100000e-08 V_low
+ 5.790000000e-08 V_low
+ 5.790100000e-08 V_hig
+ 5.800000000e-08 V_hig
+ 5.800100000e-08 V_hig
+ 5.810000000e-08 V_hig
+ 5.810100000e-08 V_hig
+ 5.820000000e-08 V_hig
+ 5.820100000e-08 V_hig
+ 5.830000000e-08 V_hig
+ 5.830100000e-08 V_hig
+ 5.840000000e-08 V_hig
+ 5.840100000e-08 V_hig
+ 5.850000000e-08 V_hig
+ 5.850100000e-08 V_hig
+ 5.860000000e-08 V_hig
+ 5.860100000e-08 V_hig
+ 5.870000000e-08 V_hig
+ 5.870100000e-08 V_hig
+ 5.880000000e-08 V_hig
+ 5.880100000e-08 V_hig
+ 5.890000000e-08 V_hig
+ 5.890100000e-08 V_hig
+ 5.900000000e-08 V_hig
+ 5.900100000e-08 V_hig
+ 5.910000000e-08 V_hig
+ 5.910100000e-08 V_hig
+ 5.920000000e-08 V_hig
+ 5.920100000e-08 V_hig
+ 5.930000000e-08 V_hig
+ 5.930100000e-08 V_hig
+ 5.940000000e-08 V_hig
+ 5.940100000e-08 V_hig
+ 5.950000000e-08 V_hig
+ 5.950100000e-08 V_hig
+ 5.960000000e-08 V_hig
+ 5.960100000e-08 V_hig
+ 5.970000000e-08 V_hig
+ 5.970100000e-08 V_hig
+ 5.980000000e-08 V_hig
+ 5.980100000e-08 V_hig
+ 5.990000000e-08 V_hig
+ 5.990100000e-08 V_low
+ 6.000000000e-08 V_low
+ 6.000100000e-08 V_low
+ 6.010000000e-08 V_low
+ 6.010100000e-08 V_low
+ 6.020000000e-08 V_low
+ 6.020100000e-08 V_low
+ 6.030000000e-08 V_low
+ 6.030100000e-08 V_low
+ 6.040000000e-08 V_low
+ 6.040100000e-08 V_low
+ 6.050000000e-08 V_low
+ 6.050100000e-08 V_low
+ 6.060000000e-08 V_low
+ 6.060100000e-08 V_low
+ 6.070000000e-08 V_low
+ 6.070100000e-08 V_low
+ 6.080000000e-08 V_low
+ 6.080100000e-08 V_low
+ 6.090000000e-08 V_low
+ 6.090100000e-08 V_low
+ 6.100000000e-08 V_low
+ 6.100100000e-08 V_low
+ 6.110000000e-08 V_low
+ 6.110100000e-08 V_low
+ 6.120000000e-08 V_low
+ 6.120100000e-08 V_low
+ 6.130000000e-08 V_low
+ 6.130100000e-08 V_low
+ 6.140000000e-08 V_low
+ 6.140100000e-08 V_low
+ 6.150000000e-08 V_low
+ 6.150100000e-08 V_low
+ 6.160000000e-08 V_low
+ 6.160100000e-08 V_low
+ 6.170000000e-08 V_low
+ 6.170100000e-08 V_low
+ 6.180000000e-08 V_low
+ 6.180100000e-08 V_low
+ 6.190000000e-08 V_low
+ 6.190100000e-08 V_hig
+ 6.200000000e-08 V_hig
+ 6.200100000e-08 V_hig
+ 6.210000000e-08 V_hig
+ 6.210100000e-08 V_hig
+ 6.220000000e-08 V_hig
+ 6.220100000e-08 V_hig
+ 6.230000000e-08 V_hig
+ 6.230100000e-08 V_hig
+ 6.240000000e-08 V_hig
+ 6.240100000e-08 V_hig
+ 6.250000000e-08 V_hig
+ 6.250100000e-08 V_hig
+ 6.260000000e-08 V_hig
+ 6.260100000e-08 V_hig
+ 6.270000000e-08 V_hig
+ 6.270100000e-08 V_hig
+ 6.280000000e-08 V_hig
+ 6.280100000e-08 V_hig
+ 6.290000000e-08 V_hig
+ 6.290100000e-08 V_hig
+ 6.300000000e-08 V_hig
+ 6.300100000e-08 V_hig
+ 6.310000000e-08 V_hig
+ 6.310100000e-08 V_hig
+ 6.320000000e-08 V_hig
+ 6.320100000e-08 V_hig
+ 6.330000000e-08 V_hig
+ 6.330100000e-08 V_hig
+ 6.340000000e-08 V_hig
+ 6.340100000e-08 V_hig
+ 6.350000000e-08 V_hig
+ 6.350100000e-08 V_hig
+ 6.360000000e-08 V_hig
+ 6.360100000e-08 V_hig
+ 6.370000000e-08 V_hig
+ 6.370100000e-08 V_hig
+ 6.380000000e-08 V_hig
+ 6.380100000e-08 V_hig
+ 6.390000000e-08 V_hig
+ 6.390100000e-08 V_low
+ 6.400000000e-08 V_low
+ 6.400100000e-08 V_low
+ 6.410000000e-08 V_low
+ 6.410100000e-08 V_low
+ 6.420000000e-08 V_low
+ 6.420100000e-08 V_low
+ 6.430000000e-08 V_low
+ 6.430100000e-08 V_low
+ 6.440000000e-08 V_low
+ 6.440100000e-08 V_low
+ 6.450000000e-08 V_low
+ 6.450100000e-08 V_low
+ 6.460000000e-08 V_low
+ 6.460100000e-08 V_low
+ 6.470000000e-08 V_low
+ 6.470100000e-08 V_low
+ 6.480000000e-08 V_low
+ 6.480100000e-08 V_low
+ 6.490000000e-08 V_low
+ 6.490100000e-08 V_hig
+ 6.500000000e-08 V_hig
+ 6.500100000e-08 V_hig
+ 6.510000000e-08 V_hig
+ 6.510100000e-08 V_hig
+ 6.520000000e-08 V_hig
+ 6.520100000e-08 V_hig
+ 6.530000000e-08 V_hig
+ 6.530100000e-08 V_hig
+ 6.540000000e-08 V_hig
+ 6.540100000e-08 V_hig
+ 6.550000000e-08 V_hig
+ 6.550100000e-08 V_hig
+ 6.560000000e-08 V_hig
+ 6.560100000e-08 V_hig
+ 6.570000000e-08 V_hig
+ 6.570100000e-08 V_hig
+ 6.580000000e-08 V_hig
+ 6.580100000e-08 V_hig
+ 6.590000000e-08 V_hig
+ 6.590100000e-08 V_low
+ 6.600000000e-08 V_low
+ 6.600100000e-08 V_low
+ 6.610000000e-08 V_low
+ 6.610100000e-08 V_low
+ 6.620000000e-08 V_low
+ 6.620100000e-08 V_low
+ 6.630000000e-08 V_low
+ 6.630100000e-08 V_low
+ 6.640000000e-08 V_low
+ 6.640100000e-08 V_low
+ 6.650000000e-08 V_low
+ 6.650100000e-08 V_low
+ 6.660000000e-08 V_low
+ 6.660100000e-08 V_low
+ 6.670000000e-08 V_low
+ 6.670100000e-08 V_low
+ 6.680000000e-08 V_low
+ 6.680100000e-08 V_low
+ 6.690000000e-08 V_low
+ 6.690100000e-08 V_hig
+ 6.700000000e-08 V_hig
+ 6.700100000e-08 V_hig
+ 6.710000000e-08 V_hig
+ 6.710100000e-08 V_hig
+ 6.720000000e-08 V_hig
+ 6.720100000e-08 V_hig
+ 6.730000000e-08 V_hig
+ 6.730100000e-08 V_hig
+ 6.740000000e-08 V_hig
+ 6.740100000e-08 V_hig
+ 6.750000000e-08 V_hig
+ 6.750100000e-08 V_hig
+ 6.760000000e-08 V_hig
+ 6.760100000e-08 V_hig
+ 6.770000000e-08 V_hig
+ 6.770100000e-08 V_hig
+ 6.780000000e-08 V_hig
+ 6.780100000e-08 V_hig
+ 6.790000000e-08 V_hig
+ 6.790100000e-08 V_hig
+ 6.800000000e-08 V_hig
+ 6.800100000e-08 V_hig
+ 6.810000000e-08 V_hig
+ 6.810100000e-08 V_hig
+ 6.820000000e-08 V_hig
+ 6.820100000e-08 V_hig
+ 6.830000000e-08 V_hig
+ 6.830100000e-08 V_hig
+ 6.840000000e-08 V_hig
+ 6.840100000e-08 V_hig
+ 6.850000000e-08 V_hig
+ 6.850100000e-08 V_hig
+ 6.860000000e-08 V_hig
+ 6.860100000e-08 V_hig
+ 6.870000000e-08 V_hig
+ 6.870100000e-08 V_hig
+ 6.880000000e-08 V_hig
+ 6.880100000e-08 V_hig
+ 6.890000000e-08 V_hig
+ 6.890100000e-08 V_hig
+ 6.900000000e-08 V_hig
+ 6.900100000e-08 V_hig
+ 6.910000000e-08 V_hig
+ 6.910100000e-08 V_hig
+ 6.920000000e-08 V_hig
+ 6.920100000e-08 V_hig
+ 6.930000000e-08 V_hig
+ 6.930100000e-08 V_hig
+ 6.940000000e-08 V_hig
+ 6.940100000e-08 V_hig
+ 6.950000000e-08 V_hig
+ 6.950100000e-08 V_hig
+ 6.960000000e-08 V_hig
+ 6.960100000e-08 V_hig
+ 6.970000000e-08 V_hig
+ 6.970100000e-08 V_hig
+ 6.980000000e-08 V_hig
+ 6.980100000e-08 V_hig
+ 6.990000000e-08 V_hig
+ 6.990100000e-08 V_low
+ 7.000000000e-08 V_low
+ 7.000100000e-08 V_low
+ 7.010000000e-08 V_low
+ 7.010100000e-08 V_low
+ 7.020000000e-08 V_low
+ 7.020100000e-08 V_low
+ 7.030000000e-08 V_low
+ 7.030100000e-08 V_low
+ 7.040000000e-08 V_low
+ 7.040100000e-08 V_low
+ 7.050000000e-08 V_low
+ 7.050100000e-08 V_low
+ 7.060000000e-08 V_low
+ 7.060100000e-08 V_low
+ 7.070000000e-08 V_low
+ 7.070100000e-08 V_low
+ 7.080000000e-08 V_low
+ 7.080100000e-08 V_low
+ 7.090000000e-08 V_low
+ 7.090100000e-08 V_low
+ 7.100000000e-08 V_low
+ 7.100100000e-08 V_low
+ 7.110000000e-08 V_low
+ 7.110100000e-08 V_low
+ 7.120000000e-08 V_low
+ 7.120100000e-08 V_low
+ 7.130000000e-08 V_low
+ 7.130100000e-08 V_low
+ 7.140000000e-08 V_low
+ 7.140100000e-08 V_low
+ 7.150000000e-08 V_low
+ 7.150100000e-08 V_low
+ 7.160000000e-08 V_low
+ 7.160100000e-08 V_low
+ 7.170000000e-08 V_low
+ 7.170100000e-08 V_low
+ 7.180000000e-08 V_low
+ 7.180100000e-08 V_low
+ 7.190000000e-08 V_low
+ 7.190100000e-08 V_hig
+ 7.200000000e-08 V_hig
+ 7.200100000e-08 V_hig
+ 7.210000000e-08 V_hig
+ 7.210100000e-08 V_hig
+ 7.220000000e-08 V_hig
+ 7.220100000e-08 V_hig
+ 7.230000000e-08 V_hig
+ 7.230100000e-08 V_hig
+ 7.240000000e-08 V_hig
+ 7.240100000e-08 V_hig
+ 7.250000000e-08 V_hig
+ 7.250100000e-08 V_hig
+ 7.260000000e-08 V_hig
+ 7.260100000e-08 V_hig
+ 7.270000000e-08 V_hig
+ 7.270100000e-08 V_hig
+ 7.280000000e-08 V_hig
+ 7.280100000e-08 V_hig
+ 7.290000000e-08 V_hig
+ 7.290100000e-08 V_low
+ 7.300000000e-08 V_low
+ 7.300100000e-08 V_low
+ 7.310000000e-08 V_low
+ 7.310100000e-08 V_low
+ 7.320000000e-08 V_low
+ 7.320100000e-08 V_low
+ 7.330000000e-08 V_low
+ 7.330100000e-08 V_low
+ 7.340000000e-08 V_low
+ 7.340100000e-08 V_low
+ 7.350000000e-08 V_low
+ 7.350100000e-08 V_low
+ 7.360000000e-08 V_low
+ 7.360100000e-08 V_low
+ 7.370000000e-08 V_low
+ 7.370100000e-08 V_low
+ 7.380000000e-08 V_low
+ 7.380100000e-08 V_low
+ 7.390000000e-08 V_low
+ 7.390100000e-08 V_low
+ 7.400000000e-08 V_low
+ 7.400100000e-08 V_low
+ 7.410000000e-08 V_low
+ 7.410100000e-08 V_low
+ 7.420000000e-08 V_low
+ 7.420100000e-08 V_low
+ 7.430000000e-08 V_low
+ 7.430100000e-08 V_low
+ 7.440000000e-08 V_low
+ 7.440100000e-08 V_low
+ 7.450000000e-08 V_low
+ 7.450100000e-08 V_low
+ 7.460000000e-08 V_low
+ 7.460100000e-08 V_low
+ 7.470000000e-08 V_low
+ 7.470100000e-08 V_low
+ 7.480000000e-08 V_low
+ 7.480100000e-08 V_low
+ 7.490000000e-08 V_low
+ 7.490100000e-08 V_hig
+ 7.500000000e-08 V_hig
+ 7.500100000e-08 V_hig
+ 7.510000000e-08 V_hig
+ 7.510100000e-08 V_hig
+ 7.520000000e-08 V_hig
+ 7.520100000e-08 V_hig
+ 7.530000000e-08 V_hig
+ 7.530100000e-08 V_hig
+ 7.540000000e-08 V_hig
+ 7.540100000e-08 V_hig
+ 7.550000000e-08 V_hig
+ 7.550100000e-08 V_hig
+ 7.560000000e-08 V_hig
+ 7.560100000e-08 V_hig
+ 7.570000000e-08 V_hig
+ 7.570100000e-08 V_hig
+ 7.580000000e-08 V_hig
+ 7.580100000e-08 V_hig
+ 7.590000000e-08 V_hig
+ 7.590100000e-08 V_hig
+ 7.600000000e-08 V_hig
+ 7.600100000e-08 V_hig
+ 7.610000000e-08 V_hig
+ 7.610100000e-08 V_hig
+ 7.620000000e-08 V_hig
+ 7.620100000e-08 V_hig
+ 7.630000000e-08 V_hig
+ 7.630100000e-08 V_hig
+ 7.640000000e-08 V_hig
+ 7.640100000e-08 V_hig
+ 7.650000000e-08 V_hig
+ 7.650100000e-08 V_hig
+ 7.660000000e-08 V_hig
+ 7.660100000e-08 V_hig
+ 7.670000000e-08 V_hig
+ 7.670100000e-08 V_hig
+ 7.680000000e-08 V_hig
+ 7.680100000e-08 V_hig
+ 7.690000000e-08 V_hig
+ 7.690100000e-08 V_hig
+ 7.700000000e-08 V_hig
+ 7.700100000e-08 V_hig
+ 7.710000000e-08 V_hig
+ 7.710100000e-08 V_hig
+ 7.720000000e-08 V_hig
+ 7.720100000e-08 V_hig
+ 7.730000000e-08 V_hig
+ 7.730100000e-08 V_hig
+ 7.740000000e-08 V_hig
+ 7.740100000e-08 V_hig
+ 7.750000000e-08 V_hig
+ 7.750100000e-08 V_hig
+ 7.760000000e-08 V_hig
+ 7.760100000e-08 V_hig
+ 7.770000000e-08 V_hig
+ 7.770100000e-08 V_hig
+ 7.780000000e-08 V_hig
+ 7.780100000e-08 V_hig
+ 7.790000000e-08 V_hig
+ 7.790100000e-08 V_hig
+ 7.800000000e-08 V_hig
+ 7.800100000e-08 V_hig
+ 7.810000000e-08 V_hig
+ 7.810100000e-08 V_hig
+ 7.820000000e-08 V_hig
+ 7.820100000e-08 V_hig
+ 7.830000000e-08 V_hig
+ 7.830100000e-08 V_hig
+ 7.840000000e-08 V_hig
+ 7.840100000e-08 V_hig
+ 7.850000000e-08 V_hig
+ 7.850100000e-08 V_hig
+ 7.860000000e-08 V_hig
+ 7.860100000e-08 V_hig
+ 7.870000000e-08 V_hig
+ 7.870100000e-08 V_hig
+ 7.880000000e-08 V_hig
+ 7.880100000e-08 V_hig
+ 7.890000000e-08 V_hig
+ 7.890100000e-08 V_hig
+ 7.900000000e-08 V_hig
+ 7.900100000e-08 V_hig
+ 7.910000000e-08 V_hig
+ 7.910100000e-08 V_hig
+ 7.920000000e-08 V_hig
+ 7.920100000e-08 V_hig
+ 7.930000000e-08 V_hig
+ 7.930100000e-08 V_hig
+ 7.940000000e-08 V_hig
+ 7.940100000e-08 V_hig
+ 7.950000000e-08 V_hig
+ 7.950100000e-08 V_hig
+ 7.960000000e-08 V_hig
+ 7.960100000e-08 V_hig
+ 7.970000000e-08 V_hig
+ 7.970100000e-08 V_hig
+ 7.980000000e-08 V_hig
+ 7.980100000e-08 V_hig
+ 7.990000000e-08 V_hig
+ 7.990100000e-08 V_low
+ 8.000000000e-08 V_low
+ 8.000100000e-08 V_low
+ 8.010000000e-08 V_low
+ 8.010100000e-08 V_low
+ 8.020000000e-08 V_low
+ 8.020100000e-08 V_low
+ 8.030000000e-08 V_low
+ 8.030100000e-08 V_low
+ 8.040000000e-08 V_low
+ 8.040100000e-08 V_low
+ 8.050000000e-08 V_low
+ 8.050100000e-08 V_low
+ 8.060000000e-08 V_low
+ 8.060100000e-08 V_low
+ 8.070000000e-08 V_low
+ 8.070100000e-08 V_low
+ 8.080000000e-08 V_low
+ 8.080100000e-08 V_low
+ 8.090000000e-08 V_low
+ 8.090100000e-08 V_low
+ 8.100000000e-08 V_low
+ 8.100100000e-08 V_low
+ 8.110000000e-08 V_low
+ 8.110100000e-08 V_low
+ 8.120000000e-08 V_low
+ 8.120100000e-08 V_low
+ 8.130000000e-08 V_low
+ 8.130100000e-08 V_low
+ 8.140000000e-08 V_low
+ 8.140100000e-08 V_low
+ 8.150000000e-08 V_low
+ 8.150100000e-08 V_low
+ 8.160000000e-08 V_low
+ 8.160100000e-08 V_low
+ 8.170000000e-08 V_low
+ 8.170100000e-08 V_low
+ 8.180000000e-08 V_low
+ 8.180100000e-08 V_low
+ 8.190000000e-08 V_low
+ 8.190100000e-08 V_hig
+ 8.200000000e-08 V_hig
+ 8.200100000e-08 V_hig
+ 8.210000000e-08 V_hig
+ 8.210100000e-08 V_hig
+ 8.220000000e-08 V_hig
+ 8.220100000e-08 V_hig
+ 8.230000000e-08 V_hig
+ 8.230100000e-08 V_hig
+ 8.240000000e-08 V_hig
+ 8.240100000e-08 V_hig
+ 8.250000000e-08 V_hig
+ 8.250100000e-08 V_hig
+ 8.260000000e-08 V_hig
+ 8.260100000e-08 V_hig
+ 8.270000000e-08 V_hig
+ 8.270100000e-08 V_hig
+ 8.280000000e-08 V_hig
+ 8.280100000e-08 V_hig
+ 8.290000000e-08 V_hig
+ 8.290100000e-08 V_hig
+ 8.300000000e-08 V_hig
+ 8.300100000e-08 V_hig
+ 8.310000000e-08 V_hig
+ 8.310100000e-08 V_hig
+ 8.320000000e-08 V_hig
+ 8.320100000e-08 V_hig
+ 8.330000000e-08 V_hig
+ 8.330100000e-08 V_hig
+ 8.340000000e-08 V_hig
+ 8.340100000e-08 V_hig
+ 8.350000000e-08 V_hig
+ 8.350100000e-08 V_hig
+ 8.360000000e-08 V_hig
+ 8.360100000e-08 V_hig
+ 8.370000000e-08 V_hig
+ 8.370100000e-08 V_hig
+ 8.380000000e-08 V_hig
+ 8.380100000e-08 V_hig
+ 8.390000000e-08 V_hig
+ 8.390100000e-08 V_hig
+ 8.400000000e-08 V_hig
+ 8.400100000e-08 V_hig
+ 8.410000000e-08 V_hig
+ 8.410100000e-08 V_hig
+ 8.420000000e-08 V_hig
+ 8.420100000e-08 V_hig
+ 8.430000000e-08 V_hig
+ 8.430100000e-08 V_hig
+ 8.440000000e-08 V_hig
+ 8.440100000e-08 V_hig
+ 8.450000000e-08 V_hig
+ 8.450100000e-08 V_hig
+ 8.460000000e-08 V_hig
+ 8.460100000e-08 V_hig
+ 8.470000000e-08 V_hig
+ 8.470100000e-08 V_hig
+ 8.480000000e-08 V_hig
+ 8.480100000e-08 V_hig
+ 8.490000000e-08 V_hig
+ 8.490100000e-08 V_hig
+ 8.500000000e-08 V_hig
+ 8.500100000e-08 V_hig
+ 8.510000000e-08 V_hig
+ 8.510100000e-08 V_hig
+ 8.520000000e-08 V_hig
+ 8.520100000e-08 V_hig
+ 8.530000000e-08 V_hig
+ 8.530100000e-08 V_hig
+ 8.540000000e-08 V_hig
+ 8.540100000e-08 V_hig
+ 8.550000000e-08 V_hig
+ 8.550100000e-08 V_hig
+ 8.560000000e-08 V_hig
+ 8.560100000e-08 V_hig
+ 8.570000000e-08 V_hig
+ 8.570100000e-08 V_hig
+ 8.580000000e-08 V_hig
+ 8.580100000e-08 V_hig
+ 8.590000000e-08 V_hig
+ 8.590100000e-08 V_hig
+ 8.600000000e-08 V_hig
+ 8.600100000e-08 V_hig
+ 8.610000000e-08 V_hig
+ 8.610100000e-08 V_hig
+ 8.620000000e-08 V_hig
+ 8.620100000e-08 V_hig
+ 8.630000000e-08 V_hig
+ 8.630100000e-08 V_hig
+ 8.640000000e-08 V_hig
+ 8.640100000e-08 V_hig
+ 8.650000000e-08 V_hig
+ 8.650100000e-08 V_hig
+ 8.660000000e-08 V_hig
+ 8.660100000e-08 V_hig
+ 8.670000000e-08 V_hig
+ 8.670100000e-08 V_hig
+ 8.680000000e-08 V_hig
+ 8.680100000e-08 V_hig
+ 8.690000000e-08 V_hig
+ 8.690100000e-08 V_low
+ 8.700000000e-08 V_low
+ 8.700100000e-08 V_low
+ 8.710000000e-08 V_low
+ 8.710100000e-08 V_low
+ 8.720000000e-08 V_low
+ 8.720100000e-08 V_low
+ 8.730000000e-08 V_low
+ 8.730100000e-08 V_low
+ 8.740000000e-08 V_low
+ 8.740100000e-08 V_low
+ 8.750000000e-08 V_low
+ 8.750100000e-08 V_low
+ 8.760000000e-08 V_low
+ 8.760100000e-08 V_low
+ 8.770000000e-08 V_low
+ 8.770100000e-08 V_low
+ 8.780000000e-08 V_low
+ 8.780100000e-08 V_low
+ 8.790000000e-08 V_low
+ 8.790100000e-08 V_hig
+ 8.800000000e-08 V_hig
+ 8.800100000e-08 V_hig
+ 8.810000000e-08 V_hig
+ 8.810100000e-08 V_hig
+ 8.820000000e-08 V_hig
+ 8.820100000e-08 V_hig
+ 8.830000000e-08 V_hig
+ 8.830100000e-08 V_hig
+ 8.840000000e-08 V_hig
+ 8.840100000e-08 V_hig
+ 8.850000000e-08 V_hig
+ 8.850100000e-08 V_hig
+ 8.860000000e-08 V_hig
+ 8.860100000e-08 V_hig
+ 8.870000000e-08 V_hig
+ 8.870100000e-08 V_hig
+ 8.880000000e-08 V_hig
+ 8.880100000e-08 V_hig
+ 8.890000000e-08 V_hig
+ 8.890100000e-08 V_low
+ 8.900000000e-08 V_low
+ 8.900100000e-08 V_low
+ 8.910000000e-08 V_low
+ 8.910100000e-08 V_low
+ 8.920000000e-08 V_low
+ 8.920100000e-08 V_low
+ 8.930000000e-08 V_low
+ 8.930100000e-08 V_low
+ 8.940000000e-08 V_low
+ 8.940100000e-08 V_low
+ 8.950000000e-08 V_low
+ 8.950100000e-08 V_low
+ 8.960000000e-08 V_low
+ 8.960100000e-08 V_low
+ 8.970000000e-08 V_low
+ 8.970100000e-08 V_low
+ 8.980000000e-08 V_low
+ 8.980100000e-08 V_low
+ 8.990000000e-08 V_low
+ 8.990100000e-08 V_hig
+ 9.000000000e-08 V_hig
+ 9.000100000e-08 V_hig
+ 9.010000000e-08 V_hig
+ 9.010100000e-08 V_hig
+ 9.020000000e-08 V_hig
+ 9.020100000e-08 V_hig
+ 9.030000000e-08 V_hig
+ 9.030100000e-08 V_hig
+ 9.040000000e-08 V_hig
+ 9.040100000e-08 V_hig
+ 9.050000000e-08 V_hig
+ 9.050100000e-08 V_hig
+ 9.060000000e-08 V_hig
+ 9.060100000e-08 V_hig
+ 9.070000000e-08 V_hig
+ 9.070100000e-08 V_hig
+ 9.080000000e-08 V_hig
+ 9.080100000e-08 V_hig
+ 9.090000000e-08 V_hig
+ 9.090100000e-08 V_hig
+ 9.100000000e-08 V_hig
+ 9.100100000e-08 V_hig
+ 9.110000000e-08 V_hig
+ 9.110100000e-08 V_hig
+ 9.120000000e-08 V_hig
+ 9.120100000e-08 V_hig
+ 9.130000000e-08 V_hig
+ 9.130100000e-08 V_hig
+ 9.140000000e-08 V_hig
+ 9.140100000e-08 V_hig
+ 9.150000000e-08 V_hig
+ 9.150100000e-08 V_hig
+ 9.160000000e-08 V_hig
+ 9.160100000e-08 V_hig
+ 9.170000000e-08 V_hig
+ 9.170100000e-08 V_hig
+ 9.180000000e-08 V_hig
+ 9.180100000e-08 V_hig
+ 9.190000000e-08 V_hig
+ 9.190100000e-08 V_hig
+ 9.200000000e-08 V_hig
+ 9.200100000e-08 V_hig
+ 9.210000000e-08 V_hig
+ 9.210100000e-08 V_hig
+ 9.220000000e-08 V_hig
+ 9.220100000e-08 V_hig
+ 9.230000000e-08 V_hig
+ 9.230100000e-08 V_hig
+ 9.240000000e-08 V_hig
+ 9.240100000e-08 V_hig
+ 9.250000000e-08 V_hig
+ 9.250100000e-08 V_hig
+ 9.260000000e-08 V_hig
+ 9.260100000e-08 V_hig
+ 9.270000000e-08 V_hig
+ 9.270100000e-08 V_hig
+ 9.280000000e-08 V_hig
+ 9.280100000e-08 V_hig
+ 9.290000000e-08 V_hig
+ 9.290100000e-08 V_low
+ 9.300000000e-08 V_low
+ 9.300100000e-08 V_low
+ 9.310000000e-08 V_low
+ 9.310100000e-08 V_low
+ 9.320000000e-08 V_low
+ 9.320100000e-08 V_low
+ 9.330000000e-08 V_low
+ 9.330100000e-08 V_low
+ 9.340000000e-08 V_low
+ 9.340100000e-08 V_low
+ 9.350000000e-08 V_low
+ 9.350100000e-08 V_low
+ 9.360000000e-08 V_low
+ 9.360100000e-08 V_low
+ 9.370000000e-08 V_low
+ 9.370100000e-08 V_low
+ 9.380000000e-08 V_low
+ 9.380100000e-08 V_low
+ 9.390000000e-08 V_low
+ 9.390100000e-08 V_low
+ 9.400000000e-08 V_low
+ 9.400100000e-08 V_low
+ 9.410000000e-08 V_low
+ 9.410100000e-08 V_low
+ 9.420000000e-08 V_low
+ 9.420100000e-08 V_low
+ 9.430000000e-08 V_low
+ 9.430100000e-08 V_low
+ 9.440000000e-08 V_low
+ 9.440100000e-08 V_low
+ 9.450000000e-08 V_low
+ 9.450100000e-08 V_low
+ 9.460000000e-08 V_low
+ 9.460100000e-08 V_low
+ 9.470000000e-08 V_low
+ 9.470100000e-08 V_low
+ 9.480000000e-08 V_low
+ 9.480100000e-08 V_low
+ 9.490000000e-08 V_low
+ 9.490100000e-08 V_hig
+ 9.500000000e-08 V_hig
+ 9.500100000e-08 V_hig
+ 9.510000000e-08 V_hig
+ 9.510100000e-08 V_hig
+ 9.520000000e-08 V_hig
+ 9.520100000e-08 V_hig
+ 9.530000000e-08 V_hig
+ 9.530100000e-08 V_hig
+ 9.540000000e-08 V_hig
+ 9.540100000e-08 V_hig
+ 9.550000000e-08 V_hig
+ 9.550100000e-08 V_hig
+ 9.560000000e-08 V_hig
+ 9.560100000e-08 V_hig
+ 9.570000000e-08 V_hig
+ 9.570100000e-08 V_hig
+ 9.580000000e-08 V_hig
+ 9.580100000e-08 V_hig
+ 9.590000000e-08 V_hig
+ 9.590100000e-08 V_hig
+ 9.600000000e-08 V_hig
+ 9.600100000e-08 V_hig
+ 9.610000000e-08 V_hig
+ 9.610100000e-08 V_hig
+ 9.620000000e-08 V_hig
+ 9.620100000e-08 V_hig
+ 9.630000000e-08 V_hig
+ 9.630100000e-08 V_hig
+ 9.640000000e-08 V_hig
+ 9.640100000e-08 V_hig
+ 9.650000000e-08 V_hig
+ 9.650100000e-08 V_hig
+ 9.660000000e-08 V_hig
+ 9.660100000e-08 V_hig
+ 9.670000000e-08 V_hig
+ 9.670100000e-08 V_hig
+ 9.680000000e-08 V_hig
+ 9.680100000e-08 V_hig
+ 9.690000000e-08 V_hig
+ 9.690100000e-08 V_hig
+ 9.700000000e-08 V_hig
+ 9.700100000e-08 V_hig
+ 9.710000000e-08 V_hig
+ 9.710100000e-08 V_hig
+ 9.720000000e-08 V_hig
+ 9.720100000e-08 V_hig
+ 9.730000000e-08 V_hig
+ 9.730100000e-08 V_hig
+ 9.740000000e-08 V_hig
+ 9.740100000e-08 V_hig
+ 9.750000000e-08 V_hig
+ 9.750100000e-08 V_hig
+ 9.760000000e-08 V_hig
+ 9.760100000e-08 V_hig
+ 9.770000000e-08 V_hig
+ 9.770100000e-08 V_hig
+ 9.780000000e-08 V_hig
+ 9.780100000e-08 V_hig
+ 9.790000000e-08 V_hig
+ 9.790100000e-08 V_hig
+ 9.800000000e-08 V_hig
+ 9.800100000e-08 V_hig
+ 9.810000000e-08 V_hig
+ 9.810100000e-08 V_hig
+ 9.820000000e-08 V_hig
+ 9.820100000e-08 V_hig
+ 9.830000000e-08 V_hig
+ 9.830100000e-08 V_hig
+ 9.840000000e-08 V_hig
+ 9.840100000e-08 V_hig
+ 9.850000000e-08 V_hig
+ 9.850100000e-08 V_hig
+ 9.860000000e-08 V_hig
+ 9.860100000e-08 V_hig
+ 9.870000000e-08 V_hig
+ 9.870100000e-08 V_hig
+ 9.880000000e-08 V_hig
+ 9.880100000e-08 V_hig
+ 9.890000000e-08 V_hig
+ 9.890100000e-08 V_low
+ 9.900000000e-08 V_low
+ 9.900100000e-08 V_low
+ 9.910000000e-08 V_low
+ 9.910100000e-08 V_low
+ 9.920000000e-08 V_low
+ 9.920100000e-08 V_low
+ 9.930000000e-08 V_low
+ 9.930100000e-08 V_low
+ 9.940000000e-08 V_low
+ 9.940100000e-08 V_low
+ 9.950000000e-08 V_low
+ 9.950100000e-08 V_low
+ 9.960000000e-08 V_low
+ 9.960100000e-08 V_low
+ 9.970000000e-08 V_low
+ 9.970100000e-08 V_low
+ 9.980000000e-08 V_low
+ 9.980100000e-08 V_low
+ 9.990000000e-08 V_low
+ 9.990100000e-08 V_hig
+ 1.000000000e-07 V_hig
+ 1.000010000e-07 V_hig
+ 1.001000000e-07 V_hig
+ 1.001010000e-07 V_hig
+ 1.002000000e-07 V_hig
+ 1.002010000e-07 V_hig
+ 1.003000000e-07 V_hig
+ 1.003010000e-07 V_hig
+ 1.004000000e-07 V_hig
+ 1.004010000e-07 V_hig
+ 1.005000000e-07 V_hig
+ 1.005010000e-07 V_hig
+ 1.006000000e-07 V_hig
+ 1.006010000e-07 V_hig
+ 1.007000000e-07 V_hig
+ 1.007010000e-07 V_hig
+ 1.008000000e-07 V_hig
+ 1.008010000e-07 V_hig
+ 1.009000000e-07 V_hig
+ 1.009010000e-07 V_hig
+ 1.010000000e-07 V_hig
+ 1.010010000e-07 V_hig
+ 1.011000000e-07 V_hig
+ 1.011010000e-07 V_hig
+ 1.012000000e-07 V_hig
+ 1.012010000e-07 V_hig
+ 1.013000000e-07 V_hig
+ 1.013010000e-07 V_hig
+ 1.014000000e-07 V_hig
+ 1.014010000e-07 V_hig
+ 1.015000000e-07 V_hig
+ 1.015010000e-07 V_hig
+ 1.016000000e-07 V_hig
+ 1.016010000e-07 V_hig
+ 1.017000000e-07 V_hig
+ 1.017010000e-07 V_hig
+ 1.018000000e-07 V_hig
+ 1.018010000e-07 V_hig
+ 1.019000000e-07 V_hig
+ 1.019010000e-07 V_low
+ 1.020000000e-07 V_low
+ 1.020010000e-07 V_low
+ 1.021000000e-07 V_low
+ 1.021010000e-07 V_low
+ 1.022000000e-07 V_low
+ 1.022010000e-07 V_low
+ 1.023000000e-07 V_low
+ 1.023010000e-07 V_low
+ 1.024000000e-07 V_low
+ 1.024010000e-07 V_low
+ 1.025000000e-07 V_low
+ 1.025010000e-07 V_low
+ 1.026000000e-07 V_low
+ 1.026010000e-07 V_low
+ 1.027000000e-07 V_low
+ 1.027010000e-07 V_low
+ 1.028000000e-07 V_low
+ 1.028010000e-07 V_low
+ 1.029000000e-07 V_low
+ 1.029010000e-07 V_low
+ 1.030000000e-07 V_low
+ 1.030010000e-07 V_low
+ 1.031000000e-07 V_low
+ 1.031010000e-07 V_low
+ 1.032000000e-07 V_low
+ 1.032010000e-07 V_low
+ 1.033000000e-07 V_low
+ 1.033010000e-07 V_low
+ 1.034000000e-07 V_low
+ 1.034010000e-07 V_low
+ 1.035000000e-07 V_low
+ 1.035010000e-07 V_low
+ 1.036000000e-07 V_low
+ 1.036010000e-07 V_low
+ 1.037000000e-07 V_low
+ 1.037010000e-07 V_low
+ 1.038000000e-07 V_low
+ 1.038010000e-07 V_low
+ 1.039000000e-07 V_low
+ 1.039010000e-07 V_hig
+ 1.040000000e-07 V_hig
+ 1.040010000e-07 V_hig
+ 1.041000000e-07 V_hig
+ 1.041010000e-07 V_hig
+ 1.042000000e-07 V_hig
+ 1.042010000e-07 V_hig
+ 1.043000000e-07 V_hig
+ 1.043010000e-07 V_hig
+ 1.044000000e-07 V_hig
+ 1.044010000e-07 V_hig
+ 1.045000000e-07 V_hig
+ 1.045010000e-07 V_hig
+ 1.046000000e-07 V_hig
+ 1.046010000e-07 V_hig
+ 1.047000000e-07 V_hig
+ 1.047010000e-07 V_hig
+ 1.048000000e-07 V_hig
+ 1.048010000e-07 V_hig
+ 1.049000000e-07 V_hig
+ 1.049010000e-07 V_low
+ 1.050000000e-07 V_low
+ 1.050010000e-07 V_low
+ 1.051000000e-07 V_low
+ 1.051010000e-07 V_low
+ 1.052000000e-07 V_low
+ 1.052010000e-07 V_low
+ 1.053000000e-07 V_low
+ 1.053010000e-07 V_low
+ 1.054000000e-07 V_low
+ 1.054010000e-07 V_low
+ 1.055000000e-07 V_low
+ 1.055010000e-07 V_low
+ 1.056000000e-07 V_low
+ 1.056010000e-07 V_low
+ 1.057000000e-07 V_low
+ 1.057010000e-07 V_low
+ 1.058000000e-07 V_low
+ 1.058010000e-07 V_low
+ 1.059000000e-07 V_low
+ 1.059010000e-07 V_low
+ 1.060000000e-07 V_low
+ 1.060010000e-07 V_low
+ 1.061000000e-07 V_low
+ 1.061010000e-07 V_low
+ 1.062000000e-07 V_low
+ 1.062010000e-07 V_low
+ 1.063000000e-07 V_low
+ 1.063010000e-07 V_low
+ 1.064000000e-07 V_low
+ 1.064010000e-07 V_low
+ 1.065000000e-07 V_low
+ 1.065010000e-07 V_low
+ 1.066000000e-07 V_low
+ 1.066010000e-07 V_low
+ 1.067000000e-07 V_low
+ 1.067010000e-07 V_low
+ 1.068000000e-07 V_low
+ 1.068010000e-07 V_low
+ 1.069000000e-07 V_low
+ 1.069010000e-07 V_hig
+ 1.070000000e-07 V_hig
+ 1.070010000e-07 V_hig
+ 1.071000000e-07 V_hig
+ 1.071010000e-07 V_hig
+ 1.072000000e-07 V_hig
+ 1.072010000e-07 V_hig
+ 1.073000000e-07 V_hig
+ 1.073010000e-07 V_hig
+ 1.074000000e-07 V_hig
+ 1.074010000e-07 V_hig
+ 1.075000000e-07 V_hig
+ 1.075010000e-07 V_hig
+ 1.076000000e-07 V_hig
+ 1.076010000e-07 V_hig
+ 1.077000000e-07 V_hig
+ 1.077010000e-07 V_hig
+ 1.078000000e-07 V_hig
+ 1.078010000e-07 V_hig
+ 1.079000000e-07 V_hig
+ 1.079010000e-07 V_hig
+ 1.080000000e-07 V_hig
+ 1.080010000e-07 V_hig
+ 1.081000000e-07 V_hig
+ 1.081010000e-07 V_hig
+ 1.082000000e-07 V_hig
+ 1.082010000e-07 V_hig
+ 1.083000000e-07 V_hig
+ 1.083010000e-07 V_hig
+ 1.084000000e-07 V_hig
+ 1.084010000e-07 V_hig
+ 1.085000000e-07 V_hig
+ 1.085010000e-07 V_hig
+ 1.086000000e-07 V_hig
+ 1.086010000e-07 V_hig
+ 1.087000000e-07 V_hig
+ 1.087010000e-07 V_hig
+ 1.088000000e-07 V_hig
+ 1.088010000e-07 V_hig
+ 1.089000000e-07 V_hig
+ 1.089010000e-07 V_low
+ 1.090000000e-07 V_low
+ 1.090010000e-07 V_low
+ 1.091000000e-07 V_low
+ 1.091010000e-07 V_low
+ 1.092000000e-07 V_low
+ 1.092010000e-07 V_low
+ 1.093000000e-07 V_low
+ 1.093010000e-07 V_low
+ 1.094000000e-07 V_low
+ 1.094010000e-07 V_low
+ 1.095000000e-07 V_low
+ 1.095010000e-07 V_low
+ 1.096000000e-07 V_low
+ 1.096010000e-07 V_low
+ 1.097000000e-07 V_low
+ 1.097010000e-07 V_low
+ 1.098000000e-07 V_low
+ 1.098010000e-07 V_low
+ 1.099000000e-07 V_low
+ 1.099010000e-07 V_hig
+ 1.100000000e-07 V_hig
+ 1.100010000e-07 V_hig
+ 1.101000000e-07 V_hig
+ 1.101010000e-07 V_hig
+ 1.102000000e-07 V_hig
+ 1.102010000e-07 V_hig
+ 1.103000000e-07 V_hig
+ 1.103010000e-07 V_hig
+ 1.104000000e-07 V_hig
+ 1.104010000e-07 V_hig
+ 1.105000000e-07 V_hig
+ 1.105010000e-07 V_hig
+ 1.106000000e-07 V_hig
+ 1.106010000e-07 V_hig
+ 1.107000000e-07 V_hig
+ 1.107010000e-07 V_hig
+ 1.108000000e-07 V_hig
+ 1.108010000e-07 V_hig
+ 1.109000000e-07 V_hig
+ 1.109010000e-07 V_hig
+ 1.110000000e-07 V_hig
+ 1.110010000e-07 V_hig
+ 1.111000000e-07 V_hig
+ 1.111010000e-07 V_hig
+ 1.112000000e-07 V_hig
+ 1.112010000e-07 V_hig
+ 1.113000000e-07 V_hig
+ 1.113010000e-07 V_hig
+ 1.114000000e-07 V_hig
+ 1.114010000e-07 V_hig
+ 1.115000000e-07 V_hig
+ 1.115010000e-07 V_hig
+ 1.116000000e-07 V_hig
+ 1.116010000e-07 V_hig
+ 1.117000000e-07 V_hig
+ 1.117010000e-07 V_hig
+ 1.118000000e-07 V_hig
+ 1.118010000e-07 V_hig
+ 1.119000000e-07 V_hig
+ 1.119010000e-07 V_hig
+ 1.120000000e-07 V_hig
+ 1.120010000e-07 V_hig
+ 1.121000000e-07 V_hig
+ 1.121010000e-07 V_hig
+ 1.122000000e-07 V_hig
+ 1.122010000e-07 V_hig
+ 1.123000000e-07 V_hig
+ 1.123010000e-07 V_hig
+ 1.124000000e-07 V_hig
+ 1.124010000e-07 V_hig
+ 1.125000000e-07 V_hig
+ 1.125010000e-07 V_hig
+ 1.126000000e-07 V_hig
+ 1.126010000e-07 V_hig
+ 1.127000000e-07 V_hig
+ 1.127010000e-07 V_hig
+ 1.128000000e-07 V_hig
+ 1.128010000e-07 V_hig
+ 1.129000000e-07 V_hig
+ 1.129010000e-07 V_hig
+ 1.130000000e-07 V_hig
+ 1.130010000e-07 V_hig
+ 1.131000000e-07 V_hig
+ 1.131010000e-07 V_hig
+ 1.132000000e-07 V_hig
+ 1.132010000e-07 V_hig
+ 1.133000000e-07 V_hig
+ 1.133010000e-07 V_hig
+ 1.134000000e-07 V_hig
+ 1.134010000e-07 V_hig
+ 1.135000000e-07 V_hig
+ 1.135010000e-07 V_hig
+ 1.136000000e-07 V_hig
+ 1.136010000e-07 V_hig
+ 1.137000000e-07 V_hig
+ 1.137010000e-07 V_hig
+ 1.138000000e-07 V_hig
+ 1.138010000e-07 V_hig
+ 1.139000000e-07 V_hig
+ 1.139010000e-07 V_hig
+ 1.140000000e-07 V_hig
+ 1.140010000e-07 V_hig
+ 1.141000000e-07 V_hig
+ 1.141010000e-07 V_hig
+ 1.142000000e-07 V_hig
+ 1.142010000e-07 V_hig
+ 1.143000000e-07 V_hig
+ 1.143010000e-07 V_hig
+ 1.144000000e-07 V_hig
+ 1.144010000e-07 V_hig
+ 1.145000000e-07 V_hig
+ 1.145010000e-07 V_hig
+ 1.146000000e-07 V_hig
+ 1.146010000e-07 V_hig
+ 1.147000000e-07 V_hig
+ 1.147010000e-07 V_hig
+ 1.148000000e-07 V_hig
+ 1.148010000e-07 V_hig
+ 1.149000000e-07 V_hig
+ 1.149010000e-07 V_hig
+ 1.150000000e-07 V_hig
+ 1.150010000e-07 V_hig
+ 1.151000000e-07 V_hig
+ 1.151010000e-07 V_hig
+ 1.152000000e-07 V_hig
+ 1.152010000e-07 V_hig
+ 1.153000000e-07 V_hig
+ 1.153010000e-07 V_hig
+ 1.154000000e-07 V_hig
+ 1.154010000e-07 V_hig
+ 1.155000000e-07 V_hig
+ 1.155010000e-07 V_hig
+ 1.156000000e-07 V_hig
+ 1.156010000e-07 V_hig
+ 1.157000000e-07 V_hig
+ 1.157010000e-07 V_hig
+ 1.158000000e-07 V_hig
+ 1.158010000e-07 V_hig
+ 1.159000000e-07 V_hig
+ 1.159010000e-07 V_hig
+ 1.160000000e-07 V_hig
+ 1.160010000e-07 V_hig
+ 1.161000000e-07 V_hig
+ 1.161010000e-07 V_hig
+ 1.162000000e-07 V_hig
+ 1.162010000e-07 V_hig
+ 1.163000000e-07 V_hig
+ 1.163010000e-07 V_hig
+ 1.164000000e-07 V_hig
+ 1.164010000e-07 V_hig
+ 1.165000000e-07 V_hig
+ 1.165010000e-07 V_hig
+ 1.166000000e-07 V_hig
+ 1.166010000e-07 V_hig
+ 1.167000000e-07 V_hig
+ 1.167010000e-07 V_hig
+ 1.168000000e-07 V_hig
+ 1.168010000e-07 V_hig
+ 1.169000000e-07 V_hig
+ 1.169010000e-07 V_hig
+ 1.170000000e-07 V_hig
+ 1.170010000e-07 V_hig
+ 1.171000000e-07 V_hig
+ 1.171010000e-07 V_hig
+ 1.172000000e-07 V_hig
+ 1.172010000e-07 V_hig
+ 1.173000000e-07 V_hig
+ 1.173010000e-07 V_hig
+ 1.174000000e-07 V_hig
+ 1.174010000e-07 V_hig
+ 1.175000000e-07 V_hig
+ 1.175010000e-07 V_hig
+ 1.176000000e-07 V_hig
+ 1.176010000e-07 V_hig
+ 1.177000000e-07 V_hig
+ 1.177010000e-07 V_hig
+ 1.178000000e-07 V_hig
+ 1.178010000e-07 V_hig
+ 1.179000000e-07 V_hig
+ 1.179010000e-07 V_hig
+ 1.180000000e-07 V_hig
+ 1.180010000e-07 V_hig
+ 1.181000000e-07 V_hig
+ 1.181010000e-07 V_hig
+ 1.182000000e-07 V_hig
+ 1.182010000e-07 V_hig
+ 1.183000000e-07 V_hig
+ 1.183010000e-07 V_hig
+ 1.184000000e-07 V_hig
+ 1.184010000e-07 V_hig
+ 1.185000000e-07 V_hig
+ 1.185010000e-07 V_hig
+ 1.186000000e-07 V_hig
+ 1.186010000e-07 V_hig
+ 1.187000000e-07 V_hig
+ 1.187010000e-07 V_hig
+ 1.188000000e-07 V_hig
+ 1.188010000e-07 V_hig
+ 1.189000000e-07 V_hig
+ 1.189010000e-07 V_low
+ 1.190000000e-07 V_low
+ 1.190010000e-07 V_low
+ 1.191000000e-07 V_low
+ 1.191010000e-07 V_low
+ 1.192000000e-07 V_low
+ 1.192010000e-07 V_low
+ 1.193000000e-07 V_low
+ 1.193010000e-07 V_low
+ 1.194000000e-07 V_low
+ 1.194010000e-07 V_low
+ 1.195000000e-07 V_low
+ 1.195010000e-07 V_low
+ 1.196000000e-07 V_low
+ 1.196010000e-07 V_low
+ 1.197000000e-07 V_low
+ 1.197010000e-07 V_low
+ 1.198000000e-07 V_low
+ 1.198010000e-07 V_low
+ 1.199000000e-07 V_low
+ 1.199010000e-07 V_hig
+ 1.200000000e-07 V_hig
+ 1.200010000e-07 V_hig
+ 1.201000000e-07 V_hig
+ 1.201010000e-07 V_hig
+ 1.202000000e-07 V_hig
+ 1.202010000e-07 V_hig
+ 1.203000000e-07 V_hig
+ 1.203010000e-07 V_hig
+ 1.204000000e-07 V_hig
+ 1.204010000e-07 V_hig
+ 1.205000000e-07 V_hig
+ 1.205010000e-07 V_hig
+ 1.206000000e-07 V_hig
+ 1.206010000e-07 V_hig
+ 1.207000000e-07 V_hig
+ 1.207010000e-07 V_hig
+ 1.208000000e-07 V_hig
+ 1.208010000e-07 V_hig
+ 1.209000000e-07 V_hig
+ 1.209010000e-07 V_hig
+ 1.210000000e-07 V_hig
+ 1.210010000e-07 V_hig
+ 1.211000000e-07 V_hig
+ 1.211010000e-07 V_hig
+ 1.212000000e-07 V_hig
+ 1.212010000e-07 V_hig
+ 1.213000000e-07 V_hig
+ 1.213010000e-07 V_hig
+ 1.214000000e-07 V_hig
+ 1.214010000e-07 V_hig
+ 1.215000000e-07 V_hig
+ 1.215010000e-07 V_hig
+ 1.216000000e-07 V_hig
+ 1.216010000e-07 V_hig
+ 1.217000000e-07 V_hig
+ 1.217010000e-07 V_hig
+ 1.218000000e-07 V_hig
+ 1.218010000e-07 V_hig
+ 1.219000000e-07 V_hig
+ 1.219010000e-07 V_low
+ 1.220000000e-07 V_low
+ 1.220010000e-07 V_low
+ 1.221000000e-07 V_low
+ 1.221010000e-07 V_low
+ 1.222000000e-07 V_low
+ 1.222010000e-07 V_low
+ 1.223000000e-07 V_low
+ 1.223010000e-07 V_low
+ 1.224000000e-07 V_low
+ 1.224010000e-07 V_low
+ 1.225000000e-07 V_low
+ 1.225010000e-07 V_low
+ 1.226000000e-07 V_low
+ 1.226010000e-07 V_low
+ 1.227000000e-07 V_low
+ 1.227010000e-07 V_low
+ 1.228000000e-07 V_low
+ 1.228010000e-07 V_low
+ 1.229000000e-07 V_low
+ 1.229010000e-07 V_hig
+ 1.230000000e-07 V_hig
+ 1.230010000e-07 V_hig
+ 1.231000000e-07 V_hig
+ 1.231010000e-07 V_hig
+ 1.232000000e-07 V_hig
+ 1.232010000e-07 V_hig
+ 1.233000000e-07 V_hig
+ 1.233010000e-07 V_hig
+ 1.234000000e-07 V_hig
+ 1.234010000e-07 V_hig
+ 1.235000000e-07 V_hig
+ 1.235010000e-07 V_hig
+ 1.236000000e-07 V_hig
+ 1.236010000e-07 V_hig
+ 1.237000000e-07 V_hig
+ 1.237010000e-07 V_hig
+ 1.238000000e-07 V_hig
+ 1.238010000e-07 V_hig
+ 1.239000000e-07 V_hig
+ 1.239010000e-07 V_low
+ 1.240000000e-07 V_low
+ 1.240010000e-07 V_low
+ 1.241000000e-07 V_low
+ 1.241010000e-07 V_low
+ 1.242000000e-07 V_low
+ 1.242010000e-07 V_low
+ 1.243000000e-07 V_low
+ 1.243010000e-07 V_low
+ 1.244000000e-07 V_low
+ 1.244010000e-07 V_low
+ 1.245000000e-07 V_low
+ 1.245010000e-07 V_low
+ 1.246000000e-07 V_low
+ 1.246010000e-07 V_low
+ 1.247000000e-07 V_low
+ 1.247010000e-07 V_low
+ 1.248000000e-07 V_low
+ 1.248010000e-07 V_low
+ 1.249000000e-07 V_low
+ 1.249010000e-07 V_low
+ 1.250000000e-07 V_low
+ 1.250010000e-07 V_low
+ 1.251000000e-07 V_low
+ 1.251010000e-07 V_low
+ 1.252000000e-07 V_low
+ 1.252010000e-07 V_low
+ 1.253000000e-07 V_low
+ 1.253010000e-07 V_low
+ 1.254000000e-07 V_low
+ 1.254010000e-07 V_low
+ 1.255000000e-07 V_low
+ 1.255010000e-07 V_low
+ 1.256000000e-07 V_low
+ 1.256010000e-07 V_low
+ 1.257000000e-07 V_low
+ 1.257010000e-07 V_low
+ 1.258000000e-07 V_low
+ 1.258010000e-07 V_low
+ 1.259000000e-07 V_low
+ 1.259010000e-07 V_hig
+ 1.260000000e-07 V_hig
+ 1.260010000e-07 V_hig
+ 1.261000000e-07 V_hig
+ 1.261010000e-07 V_hig
+ 1.262000000e-07 V_hig
+ 1.262010000e-07 V_hig
+ 1.263000000e-07 V_hig
+ 1.263010000e-07 V_hig
+ 1.264000000e-07 V_hig
+ 1.264010000e-07 V_hig
+ 1.265000000e-07 V_hig
+ 1.265010000e-07 V_hig
+ 1.266000000e-07 V_hig
+ 1.266010000e-07 V_hig
+ 1.267000000e-07 V_hig
+ 1.267010000e-07 V_hig
+ 1.268000000e-07 V_hig
+ 1.268010000e-07 V_hig
+ 1.269000000e-07 V_hig
+ 1.269010000e-07 V_low
+ 1.270000000e-07 V_low
+ 1.270010000e-07 V_low
+ 1.271000000e-07 V_low
+ 1.271010000e-07 V_low
+ 1.272000000e-07 V_low
+ 1.272010000e-07 V_low
+ 1.273000000e-07 V_low
+ 1.273010000e-07 V_low
+ 1.274000000e-07 V_low
+ 1.274010000e-07 V_low
+ 1.275000000e-07 V_low
+ 1.275010000e-07 V_low
+ 1.276000000e-07 V_low
+ 1.276010000e-07 V_low
+ 1.277000000e-07 V_low
+ 1.277010000e-07 V_low
+ 1.278000000e-07 V_low
+ 1.278010000e-07 V_low
+ 1.279000000e-07 V_low
+ 1.279010000e-07 V_low
+ 1.280000000e-07 V_low
+ 1.280010000e-07 V_low
+ 1.281000000e-07 V_low
+ 1.281010000e-07 V_low
+ 1.282000000e-07 V_low
+ 1.282010000e-07 V_low
+ 1.283000000e-07 V_low
+ 1.283010000e-07 V_low
+ 1.284000000e-07 V_low
+ 1.284010000e-07 V_low
+ 1.285000000e-07 V_low
+ 1.285010000e-07 V_low
+ 1.286000000e-07 V_low
+ 1.286010000e-07 V_low
+ 1.287000000e-07 V_low
+ 1.287010000e-07 V_low
+ 1.288000000e-07 V_low
+ 1.288010000e-07 V_low
+ 1.289000000e-07 V_low
+ 1.289010000e-07 V_hig
+ 1.290000000e-07 V_hig
+ 1.290010000e-07 V_hig
+ 1.291000000e-07 V_hig
+ 1.291010000e-07 V_hig
+ 1.292000000e-07 V_hig
+ 1.292010000e-07 V_hig
+ 1.293000000e-07 V_hig
+ 1.293010000e-07 V_hig
+ 1.294000000e-07 V_hig
+ 1.294010000e-07 V_hig
+ 1.295000000e-07 V_hig
+ 1.295010000e-07 V_hig
+ 1.296000000e-07 V_hig
+ 1.296010000e-07 V_hig
+ 1.297000000e-07 V_hig
+ 1.297010000e-07 V_hig
+ 1.298000000e-07 V_hig
+ 1.298010000e-07 V_hig
+ 1.299000000e-07 V_hig
+ 1.299010000e-07 V_hig
+ 1.300000000e-07 V_hig
+ 1.300010000e-07 V_hig
+ 1.301000000e-07 V_hig
+ 1.301010000e-07 V_hig
+ 1.302000000e-07 V_hig
+ 1.302010000e-07 V_hig
+ 1.303000000e-07 V_hig
+ 1.303010000e-07 V_hig
+ 1.304000000e-07 V_hig
+ 1.304010000e-07 V_hig
+ 1.305000000e-07 V_hig
+ 1.305010000e-07 V_hig
+ 1.306000000e-07 V_hig
+ 1.306010000e-07 V_hig
+ 1.307000000e-07 V_hig
+ 1.307010000e-07 V_hig
+ 1.308000000e-07 V_hig
+ 1.308010000e-07 V_hig
+ 1.309000000e-07 V_hig
+ 1.309010000e-07 V_low
+ 1.310000000e-07 V_low
+ 1.310010000e-07 V_low
+ 1.311000000e-07 V_low
+ 1.311010000e-07 V_low
+ 1.312000000e-07 V_low
+ 1.312010000e-07 V_low
+ 1.313000000e-07 V_low
+ 1.313010000e-07 V_low
+ 1.314000000e-07 V_low
+ 1.314010000e-07 V_low
+ 1.315000000e-07 V_low
+ 1.315010000e-07 V_low
+ 1.316000000e-07 V_low
+ 1.316010000e-07 V_low
+ 1.317000000e-07 V_low
+ 1.317010000e-07 V_low
+ 1.318000000e-07 V_low
+ 1.318010000e-07 V_low
+ 1.319000000e-07 V_low
+ 1.319010000e-07 V_low
+ 1.320000000e-07 V_low
+ 1.320010000e-07 V_low
+ 1.321000000e-07 V_low
+ 1.321010000e-07 V_low
+ 1.322000000e-07 V_low
+ 1.322010000e-07 V_low
+ 1.323000000e-07 V_low
+ 1.323010000e-07 V_low
+ 1.324000000e-07 V_low
+ 1.324010000e-07 V_low
+ 1.325000000e-07 V_low
+ 1.325010000e-07 V_low
+ 1.326000000e-07 V_low
+ 1.326010000e-07 V_low
+ 1.327000000e-07 V_low
+ 1.327010000e-07 V_low
+ 1.328000000e-07 V_low
+ 1.328010000e-07 V_low
+ 1.329000000e-07 V_low
+ 1.329010000e-07 V_hig
+ 1.330000000e-07 V_hig
+ 1.330010000e-07 V_hig
+ 1.331000000e-07 V_hig
+ 1.331010000e-07 V_hig
+ 1.332000000e-07 V_hig
+ 1.332010000e-07 V_hig
+ 1.333000000e-07 V_hig
+ 1.333010000e-07 V_hig
+ 1.334000000e-07 V_hig
+ 1.334010000e-07 V_hig
+ 1.335000000e-07 V_hig
+ 1.335010000e-07 V_hig
+ 1.336000000e-07 V_hig
+ 1.336010000e-07 V_hig
+ 1.337000000e-07 V_hig
+ 1.337010000e-07 V_hig
+ 1.338000000e-07 V_hig
+ 1.338010000e-07 V_hig
+ 1.339000000e-07 V_hig
+ 1.339010000e-07 V_low
+ 1.340000000e-07 V_low
+ 1.340010000e-07 V_low
+ 1.341000000e-07 V_low
+ 1.341010000e-07 V_low
+ 1.342000000e-07 V_low
+ 1.342010000e-07 V_low
+ 1.343000000e-07 V_low
+ 1.343010000e-07 V_low
+ 1.344000000e-07 V_low
+ 1.344010000e-07 V_low
+ 1.345000000e-07 V_low
+ 1.345010000e-07 V_low
+ 1.346000000e-07 V_low
+ 1.346010000e-07 V_low
+ 1.347000000e-07 V_low
+ 1.347010000e-07 V_low
+ 1.348000000e-07 V_low
+ 1.348010000e-07 V_low
+ 1.349000000e-07 V_low
+ 1.349010000e-07 V_hig
+ 1.350000000e-07 V_hig
+ 1.350010000e-07 V_hig
+ 1.351000000e-07 V_hig
+ 1.351010000e-07 V_hig
+ 1.352000000e-07 V_hig
+ 1.352010000e-07 V_hig
+ 1.353000000e-07 V_hig
+ 1.353010000e-07 V_hig
+ 1.354000000e-07 V_hig
+ 1.354010000e-07 V_hig
+ 1.355000000e-07 V_hig
+ 1.355010000e-07 V_hig
+ 1.356000000e-07 V_hig
+ 1.356010000e-07 V_hig
+ 1.357000000e-07 V_hig
+ 1.357010000e-07 V_hig
+ 1.358000000e-07 V_hig
+ 1.358010000e-07 V_hig
+ 1.359000000e-07 V_hig
+ 1.359010000e-07 V_hig
+ 1.360000000e-07 V_hig
+ 1.360010000e-07 V_hig
+ 1.361000000e-07 V_hig
+ 1.361010000e-07 V_hig
+ 1.362000000e-07 V_hig
+ 1.362010000e-07 V_hig
+ 1.363000000e-07 V_hig
+ 1.363010000e-07 V_hig
+ 1.364000000e-07 V_hig
+ 1.364010000e-07 V_hig
+ 1.365000000e-07 V_hig
+ 1.365010000e-07 V_hig
+ 1.366000000e-07 V_hig
+ 1.366010000e-07 V_hig
+ 1.367000000e-07 V_hig
+ 1.367010000e-07 V_hig
+ 1.368000000e-07 V_hig
+ 1.368010000e-07 V_hig
+ 1.369000000e-07 V_hig
+ 1.369010000e-07 V_hig
+ 1.370000000e-07 V_hig
+ 1.370010000e-07 V_hig
+ 1.371000000e-07 V_hig
+ 1.371010000e-07 V_hig
+ 1.372000000e-07 V_hig
+ 1.372010000e-07 V_hig
+ 1.373000000e-07 V_hig
+ 1.373010000e-07 V_hig
+ 1.374000000e-07 V_hig
+ 1.374010000e-07 V_hig
+ 1.375000000e-07 V_hig
+ 1.375010000e-07 V_hig
+ 1.376000000e-07 V_hig
+ 1.376010000e-07 V_hig
+ 1.377000000e-07 V_hig
+ 1.377010000e-07 V_hig
+ 1.378000000e-07 V_hig
+ 1.378010000e-07 V_hig
+ 1.379000000e-07 V_hig
+ 1.379010000e-07 V_low
+ 1.380000000e-07 V_low
+ 1.380010000e-07 V_low
+ 1.381000000e-07 V_low
+ 1.381010000e-07 V_low
+ 1.382000000e-07 V_low
+ 1.382010000e-07 V_low
+ 1.383000000e-07 V_low
+ 1.383010000e-07 V_low
+ 1.384000000e-07 V_low
+ 1.384010000e-07 V_low
+ 1.385000000e-07 V_low
+ 1.385010000e-07 V_low
+ 1.386000000e-07 V_low
+ 1.386010000e-07 V_low
+ 1.387000000e-07 V_low
+ 1.387010000e-07 V_low
+ 1.388000000e-07 V_low
+ 1.388010000e-07 V_low
+ 1.389000000e-07 V_low
+ 1.389010000e-07 V_hig
+ 1.390000000e-07 V_hig
+ 1.390010000e-07 V_hig
+ 1.391000000e-07 V_hig
+ 1.391010000e-07 V_hig
+ 1.392000000e-07 V_hig
+ 1.392010000e-07 V_hig
+ 1.393000000e-07 V_hig
+ 1.393010000e-07 V_hig
+ 1.394000000e-07 V_hig
+ 1.394010000e-07 V_hig
+ 1.395000000e-07 V_hig
+ 1.395010000e-07 V_hig
+ 1.396000000e-07 V_hig
+ 1.396010000e-07 V_hig
+ 1.397000000e-07 V_hig
+ 1.397010000e-07 V_hig
+ 1.398000000e-07 V_hig
+ 1.398010000e-07 V_hig
+ 1.399000000e-07 V_hig
+ 1.399010000e-07 V_low
+ 1.400000000e-07 V_low
+ 1.400010000e-07 V_low
+ 1.401000000e-07 V_low
+ 1.401010000e-07 V_low
+ 1.402000000e-07 V_low
+ 1.402010000e-07 V_low
+ 1.403000000e-07 V_low
+ 1.403010000e-07 V_low
+ 1.404000000e-07 V_low
+ 1.404010000e-07 V_low
+ 1.405000000e-07 V_low
+ 1.405010000e-07 V_low
+ 1.406000000e-07 V_low
+ 1.406010000e-07 V_low
+ 1.407000000e-07 V_low
+ 1.407010000e-07 V_low
+ 1.408000000e-07 V_low
+ 1.408010000e-07 V_low
+ 1.409000000e-07 V_low
+ 1.409010000e-07 V_hig
+ 1.410000000e-07 V_hig
+ 1.410010000e-07 V_hig
+ 1.411000000e-07 V_hig
+ 1.411010000e-07 V_hig
+ 1.412000000e-07 V_hig
+ 1.412010000e-07 V_hig
+ 1.413000000e-07 V_hig
+ 1.413010000e-07 V_hig
+ 1.414000000e-07 V_hig
+ 1.414010000e-07 V_hig
+ 1.415000000e-07 V_hig
+ 1.415010000e-07 V_hig
+ 1.416000000e-07 V_hig
+ 1.416010000e-07 V_hig
+ 1.417000000e-07 V_hig
+ 1.417010000e-07 V_hig
+ 1.418000000e-07 V_hig
+ 1.418010000e-07 V_hig
+ 1.419000000e-07 V_hig
+ 1.419010000e-07 V_hig
+ 1.420000000e-07 V_hig
+ 1.420010000e-07 V_hig
+ 1.421000000e-07 V_hig
+ 1.421010000e-07 V_hig
+ 1.422000000e-07 V_hig
+ 1.422010000e-07 V_hig
+ 1.423000000e-07 V_hig
+ 1.423010000e-07 V_hig
+ 1.424000000e-07 V_hig
+ 1.424010000e-07 V_hig
+ 1.425000000e-07 V_hig
+ 1.425010000e-07 V_hig
+ 1.426000000e-07 V_hig
+ 1.426010000e-07 V_hig
+ 1.427000000e-07 V_hig
+ 1.427010000e-07 V_hig
+ 1.428000000e-07 V_hig
+ 1.428010000e-07 V_hig
+ 1.429000000e-07 V_hig
+ 1.429010000e-07 V_low
+ 1.430000000e-07 V_low
+ 1.430010000e-07 V_low
+ 1.431000000e-07 V_low
+ 1.431010000e-07 V_low
+ 1.432000000e-07 V_low
+ 1.432010000e-07 V_low
+ 1.433000000e-07 V_low
+ 1.433010000e-07 V_low
+ 1.434000000e-07 V_low
+ 1.434010000e-07 V_low
+ 1.435000000e-07 V_low
+ 1.435010000e-07 V_low
+ 1.436000000e-07 V_low
+ 1.436010000e-07 V_low
+ 1.437000000e-07 V_low
+ 1.437010000e-07 V_low
+ 1.438000000e-07 V_low
+ 1.438010000e-07 V_low
+ 1.439000000e-07 V_low
+ 1.439010000e-07 V_hig
+ 1.440000000e-07 V_hig
+ 1.440010000e-07 V_hig
+ 1.441000000e-07 V_hig
+ 1.441010000e-07 V_hig
+ 1.442000000e-07 V_hig
+ 1.442010000e-07 V_hig
+ 1.443000000e-07 V_hig
+ 1.443010000e-07 V_hig
+ 1.444000000e-07 V_hig
+ 1.444010000e-07 V_hig
+ 1.445000000e-07 V_hig
+ 1.445010000e-07 V_hig
+ 1.446000000e-07 V_hig
+ 1.446010000e-07 V_hig
+ 1.447000000e-07 V_hig
+ 1.447010000e-07 V_hig
+ 1.448000000e-07 V_hig
+ 1.448010000e-07 V_hig
+ 1.449000000e-07 V_hig
+ 1.449010000e-07 V_low
+ 1.450000000e-07 V_low
+ 1.450010000e-07 V_low
+ 1.451000000e-07 V_low
+ 1.451010000e-07 V_low
+ 1.452000000e-07 V_low
+ 1.452010000e-07 V_low
+ 1.453000000e-07 V_low
+ 1.453010000e-07 V_low
+ 1.454000000e-07 V_low
+ 1.454010000e-07 V_low
+ 1.455000000e-07 V_low
+ 1.455010000e-07 V_low
+ 1.456000000e-07 V_low
+ 1.456010000e-07 V_low
+ 1.457000000e-07 V_low
+ 1.457010000e-07 V_low
+ 1.458000000e-07 V_low
+ 1.458010000e-07 V_low
+ 1.459000000e-07 V_low
+ 1.459010000e-07 V_hig
+ 1.460000000e-07 V_hig
+ 1.460010000e-07 V_hig
+ 1.461000000e-07 V_hig
+ 1.461010000e-07 V_hig
+ 1.462000000e-07 V_hig
+ 1.462010000e-07 V_hig
+ 1.463000000e-07 V_hig
+ 1.463010000e-07 V_hig
+ 1.464000000e-07 V_hig
+ 1.464010000e-07 V_hig
+ 1.465000000e-07 V_hig
+ 1.465010000e-07 V_hig
+ 1.466000000e-07 V_hig
+ 1.466010000e-07 V_hig
+ 1.467000000e-07 V_hig
+ 1.467010000e-07 V_hig
+ 1.468000000e-07 V_hig
+ 1.468010000e-07 V_hig
+ 1.469000000e-07 V_hig
+ 1.469010000e-07 V_hig
+ 1.470000000e-07 V_hig
+ 1.470010000e-07 V_hig
+ 1.471000000e-07 V_hig
+ 1.471010000e-07 V_hig
+ 1.472000000e-07 V_hig
+ 1.472010000e-07 V_hig
+ 1.473000000e-07 V_hig
+ 1.473010000e-07 V_hig
+ 1.474000000e-07 V_hig
+ 1.474010000e-07 V_hig
+ 1.475000000e-07 V_hig
+ 1.475010000e-07 V_hig
+ 1.476000000e-07 V_hig
+ 1.476010000e-07 V_hig
+ 1.477000000e-07 V_hig
+ 1.477010000e-07 V_hig
+ 1.478000000e-07 V_hig
+ 1.478010000e-07 V_hig
+ 1.479000000e-07 V_hig
+ 1.479010000e-07 V_low
+ 1.480000000e-07 V_low
+ 1.480010000e-07 V_low
+ 1.481000000e-07 V_low
+ 1.481010000e-07 V_low
+ 1.482000000e-07 V_low
+ 1.482010000e-07 V_low
+ 1.483000000e-07 V_low
+ 1.483010000e-07 V_low
+ 1.484000000e-07 V_low
+ 1.484010000e-07 V_low
+ 1.485000000e-07 V_low
+ 1.485010000e-07 V_low
+ 1.486000000e-07 V_low
+ 1.486010000e-07 V_low
+ 1.487000000e-07 V_low
+ 1.487010000e-07 V_low
+ 1.488000000e-07 V_low
+ 1.488010000e-07 V_low
+ 1.489000000e-07 V_low
+ 1.489010000e-07 V_low
+ 1.490000000e-07 V_low
+ 1.490010000e-07 V_low
+ 1.491000000e-07 V_low
+ 1.491010000e-07 V_low
+ 1.492000000e-07 V_low
+ 1.492010000e-07 V_low
+ 1.493000000e-07 V_low
+ 1.493010000e-07 V_low
+ 1.494000000e-07 V_low
+ 1.494010000e-07 V_low
+ 1.495000000e-07 V_low
+ 1.495010000e-07 V_low
+ 1.496000000e-07 V_low
+ 1.496010000e-07 V_low
+ 1.497000000e-07 V_low
+ 1.497010000e-07 V_low
+ 1.498000000e-07 V_low
+ 1.498010000e-07 V_low
+ 1.499000000e-07 V_low
+ 1.499010000e-07 V_hig
+ 1.500000000e-07 V_hig
+ 1.500010000e-07 V_hig
+ 1.501000000e-07 V_hig
+ 1.501010000e-07 V_hig
+ 1.502000000e-07 V_hig
+ 1.502010000e-07 V_hig
+ 1.503000000e-07 V_hig
+ 1.503010000e-07 V_hig
+ 1.504000000e-07 V_hig
+ 1.504010000e-07 V_hig
+ 1.505000000e-07 V_hig
+ 1.505010000e-07 V_hig
+ 1.506000000e-07 V_hig
+ 1.506010000e-07 V_hig
+ 1.507000000e-07 V_hig
+ 1.507010000e-07 V_hig
+ 1.508000000e-07 V_hig
+ 1.508010000e-07 V_hig
+ 1.509000000e-07 V_hig
+ 1.509010000e-07 V_low
+ 1.510000000e-07 V_low
+ 1.510010000e-07 V_low
+ 1.511000000e-07 V_low
+ 1.511010000e-07 V_low
+ 1.512000000e-07 V_low
+ 1.512010000e-07 V_low
+ 1.513000000e-07 V_low
+ 1.513010000e-07 V_low
+ 1.514000000e-07 V_low
+ 1.514010000e-07 V_low
+ 1.515000000e-07 V_low
+ 1.515010000e-07 V_low
+ 1.516000000e-07 V_low
+ 1.516010000e-07 V_low
+ 1.517000000e-07 V_low
+ 1.517010000e-07 V_low
+ 1.518000000e-07 V_low
+ 1.518010000e-07 V_low
+ 1.519000000e-07 V_low
+ 1.519010000e-07 V_low
+ 1.520000000e-07 V_low
+ 1.520010000e-07 V_low
+ 1.521000000e-07 V_low
+ 1.521010000e-07 V_low
+ 1.522000000e-07 V_low
+ 1.522010000e-07 V_low
+ 1.523000000e-07 V_low
+ 1.523010000e-07 V_low
+ 1.524000000e-07 V_low
+ 1.524010000e-07 V_low
+ 1.525000000e-07 V_low
+ 1.525010000e-07 V_low
+ 1.526000000e-07 V_low
+ 1.526010000e-07 V_low
+ 1.527000000e-07 V_low
+ 1.527010000e-07 V_low
+ 1.528000000e-07 V_low
+ 1.528010000e-07 V_low
+ 1.529000000e-07 V_low
+ 1.529010000e-07 V_hig
+ 1.530000000e-07 V_hig
+ 1.530010000e-07 V_hig
+ 1.531000000e-07 V_hig
+ 1.531010000e-07 V_hig
+ 1.532000000e-07 V_hig
+ 1.532010000e-07 V_hig
+ 1.533000000e-07 V_hig
+ 1.533010000e-07 V_hig
+ 1.534000000e-07 V_hig
+ 1.534010000e-07 V_hig
+ 1.535000000e-07 V_hig
+ 1.535010000e-07 V_hig
+ 1.536000000e-07 V_hig
+ 1.536010000e-07 V_hig
+ 1.537000000e-07 V_hig
+ 1.537010000e-07 V_hig
+ 1.538000000e-07 V_hig
+ 1.538010000e-07 V_hig
+ 1.539000000e-07 V_hig
+ 1.539010000e-07 V_low
+ 1.540000000e-07 V_low
+ 1.540010000e-07 V_low
+ 1.541000000e-07 V_low
+ 1.541010000e-07 V_low
+ 1.542000000e-07 V_low
+ 1.542010000e-07 V_low
+ 1.543000000e-07 V_low
+ 1.543010000e-07 V_low
+ 1.544000000e-07 V_low
+ 1.544010000e-07 V_low
+ 1.545000000e-07 V_low
+ 1.545010000e-07 V_low
+ 1.546000000e-07 V_low
+ 1.546010000e-07 V_low
+ 1.547000000e-07 V_low
+ 1.547010000e-07 V_low
+ 1.548000000e-07 V_low
+ 1.548010000e-07 V_low
+ 1.549000000e-07 V_low
+ 1.549010000e-07 V_low
+ 1.550000000e-07 V_low
+ 1.550010000e-07 V_low
+ 1.551000000e-07 V_low
+ 1.551010000e-07 V_low
+ 1.552000000e-07 V_low
+ 1.552010000e-07 V_low
+ 1.553000000e-07 V_low
+ 1.553010000e-07 V_low
+ 1.554000000e-07 V_low
+ 1.554010000e-07 V_low
+ 1.555000000e-07 V_low
+ 1.555010000e-07 V_low
+ 1.556000000e-07 V_low
+ 1.556010000e-07 V_low
+ 1.557000000e-07 V_low
+ 1.557010000e-07 V_low
+ 1.558000000e-07 V_low
+ 1.558010000e-07 V_low
+ 1.559000000e-07 V_low
+ 1.559010000e-07 V_low
+ 1.560000000e-07 V_low
+ 1.560010000e-07 V_low
+ 1.561000000e-07 V_low
+ 1.561010000e-07 V_low
+ 1.562000000e-07 V_low
+ 1.562010000e-07 V_low
+ 1.563000000e-07 V_low
+ 1.563010000e-07 V_low
+ 1.564000000e-07 V_low
+ 1.564010000e-07 V_low
+ 1.565000000e-07 V_low
+ 1.565010000e-07 V_low
+ 1.566000000e-07 V_low
+ 1.566010000e-07 V_low
+ 1.567000000e-07 V_low
+ 1.567010000e-07 V_low
+ 1.568000000e-07 V_low
+ 1.568010000e-07 V_low
+ 1.569000000e-07 V_low
+ 1.569010000e-07 V_hig
+ 1.570000000e-07 V_hig
+ 1.570010000e-07 V_hig
+ 1.571000000e-07 V_hig
+ 1.571010000e-07 V_hig
+ 1.572000000e-07 V_hig
+ 1.572010000e-07 V_hig
+ 1.573000000e-07 V_hig
+ 1.573010000e-07 V_hig
+ 1.574000000e-07 V_hig
+ 1.574010000e-07 V_hig
+ 1.575000000e-07 V_hig
+ 1.575010000e-07 V_hig
+ 1.576000000e-07 V_hig
+ 1.576010000e-07 V_hig
+ 1.577000000e-07 V_hig
+ 1.577010000e-07 V_hig
+ 1.578000000e-07 V_hig
+ 1.578010000e-07 V_hig
+ 1.579000000e-07 V_hig
+ 1.579010000e-07 V_low
+ 1.580000000e-07 V_low
+ 1.580010000e-07 V_low
+ 1.581000000e-07 V_low
+ 1.581010000e-07 V_low
+ 1.582000000e-07 V_low
+ 1.582010000e-07 V_low
+ 1.583000000e-07 V_low
+ 1.583010000e-07 V_low
+ 1.584000000e-07 V_low
+ 1.584010000e-07 V_low
+ 1.585000000e-07 V_low
+ 1.585010000e-07 V_low
+ 1.586000000e-07 V_low
+ 1.586010000e-07 V_low
+ 1.587000000e-07 V_low
+ 1.587010000e-07 V_low
+ 1.588000000e-07 V_low
+ 1.588010000e-07 V_low
+ 1.589000000e-07 V_low
+ 1.589010000e-07 V_low
+ 1.590000000e-07 V_low
+ 1.590010000e-07 V_low
+ 1.591000000e-07 V_low
+ 1.591010000e-07 V_low
+ 1.592000000e-07 V_low
+ 1.592010000e-07 V_low
+ 1.593000000e-07 V_low
+ 1.593010000e-07 V_low
+ 1.594000000e-07 V_low
+ 1.594010000e-07 V_low
+ 1.595000000e-07 V_low
+ 1.595010000e-07 V_low
+ 1.596000000e-07 V_low
+ 1.596010000e-07 V_low
+ 1.597000000e-07 V_low
+ 1.597010000e-07 V_low
+ 1.598000000e-07 V_low
+ 1.598010000e-07 V_low
+ 1.599000000e-07 V_low
+ 1.599010000e-07 V_hig
+ 1.600000000e-07 V_hig
+ 1.600010000e-07 V_hig
+ 1.601000000e-07 V_hig
+ 1.601010000e-07 V_hig
+ 1.602000000e-07 V_hig
+ 1.602010000e-07 V_hig
+ 1.603000000e-07 V_hig
+ 1.603010000e-07 V_hig
+ 1.604000000e-07 V_hig
+ 1.604010000e-07 V_hig
+ 1.605000000e-07 V_hig
+ 1.605010000e-07 V_hig
+ 1.606000000e-07 V_hig
+ 1.606010000e-07 V_hig
+ 1.607000000e-07 V_hig
+ 1.607010000e-07 V_hig
+ 1.608000000e-07 V_hig
+ 1.608010000e-07 V_hig
+ 1.609000000e-07 V_hig
+ 1.609010000e-07 V_low
+ 1.610000000e-07 V_low
+ 1.610010000e-07 V_low
+ 1.611000000e-07 V_low
+ 1.611010000e-07 V_low
+ 1.612000000e-07 V_low
+ 1.612010000e-07 V_low
+ 1.613000000e-07 V_low
+ 1.613010000e-07 V_low
+ 1.614000000e-07 V_low
+ 1.614010000e-07 V_low
+ 1.615000000e-07 V_low
+ 1.615010000e-07 V_low
+ 1.616000000e-07 V_low
+ 1.616010000e-07 V_low
+ 1.617000000e-07 V_low
+ 1.617010000e-07 V_low
+ 1.618000000e-07 V_low
+ 1.618010000e-07 V_low
+ 1.619000000e-07 V_low
+ 1.619010000e-07 V_low
+ 1.620000000e-07 V_low
+ 1.620010000e-07 V_low
+ 1.621000000e-07 V_low
+ 1.621010000e-07 V_low
+ 1.622000000e-07 V_low
+ 1.622010000e-07 V_low
+ 1.623000000e-07 V_low
+ 1.623010000e-07 V_low
+ 1.624000000e-07 V_low
+ 1.624010000e-07 V_low
+ 1.625000000e-07 V_low
+ 1.625010000e-07 V_low
+ 1.626000000e-07 V_low
+ 1.626010000e-07 V_low
+ 1.627000000e-07 V_low
+ 1.627010000e-07 V_low
+ 1.628000000e-07 V_low
+ 1.628010000e-07 V_low
+ 1.629000000e-07 V_low
+ 1.629010000e-07 V_hig
+ 1.630000000e-07 V_hig
+ 1.630010000e-07 V_hig
+ 1.631000000e-07 V_hig
+ 1.631010000e-07 V_hig
+ 1.632000000e-07 V_hig
+ 1.632010000e-07 V_hig
+ 1.633000000e-07 V_hig
+ 1.633010000e-07 V_hig
+ 1.634000000e-07 V_hig
+ 1.634010000e-07 V_hig
+ 1.635000000e-07 V_hig
+ 1.635010000e-07 V_hig
+ 1.636000000e-07 V_hig
+ 1.636010000e-07 V_hig
+ 1.637000000e-07 V_hig
+ 1.637010000e-07 V_hig
+ 1.638000000e-07 V_hig
+ 1.638010000e-07 V_hig
+ 1.639000000e-07 V_hig
+ 1.639010000e-07 V_low
+ 1.640000000e-07 V_low
+ 1.640010000e-07 V_low
+ 1.641000000e-07 V_low
+ 1.641010000e-07 V_low
+ 1.642000000e-07 V_low
+ 1.642010000e-07 V_low
+ 1.643000000e-07 V_low
+ 1.643010000e-07 V_low
+ 1.644000000e-07 V_low
+ 1.644010000e-07 V_low
+ 1.645000000e-07 V_low
+ 1.645010000e-07 V_low
+ 1.646000000e-07 V_low
+ 1.646010000e-07 V_low
+ 1.647000000e-07 V_low
+ 1.647010000e-07 V_low
+ 1.648000000e-07 V_low
+ 1.648010000e-07 V_low
+ 1.649000000e-07 V_low
+ 1.649010000e-07 V_low
+ 1.650000000e-07 V_low
+ 1.650010000e-07 V_low
+ 1.651000000e-07 V_low
+ 1.651010000e-07 V_low
+ 1.652000000e-07 V_low
+ 1.652010000e-07 V_low
+ 1.653000000e-07 V_low
+ 1.653010000e-07 V_low
+ 1.654000000e-07 V_low
+ 1.654010000e-07 V_low
+ 1.655000000e-07 V_low
+ 1.655010000e-07 V_low
+ 1.656000000e-07 V_low
+ 1.656010000e-07 V_low
+ 1.657000000e-07 V_low
+ 1.657010000e-07 V_low
+ 1.658000000e-07 V_low
+ 1.658010000e-07 V_low
+ 1.659000000e-07 V_low
+ 1.659010000e-07 V_low
+ 1.660000000e-07 V_low
+ 1.660010000e-07 V_low
+ 1.661000000e-07 V_low
+ 1.661010000e-07 V_low
+ 1.662000000e-07 V_low
+ 1.662010000e-07 V_low
+ 1.663000000e-07 V_low
+ 1.663010000e-07 V_low
+ 1.664000000e-07 V_low
+ 1.664010000e-07 V_low
+ 1.665000000e-07 V_low
+ 1.665010000e-07 V_low
+ 1.666000000e-07 V_low
+ 1.666010000e-07 V_low
+ 1.667000000e-07 V_low
+ 1.667010000e-07 V_low
+ 1.668000000e-07 V_low
+ 1.668010000e-07 V_low
+ 1.669000000e-07 V_low
+ 1.669010000e-07 V_low
+ 1.670000000e-07 V_low
+ 1.670010000e-07 V_low
+ 1.671000000e-07 V_low
+ 1.671010000e-07 V_low
+ 1.672000000e-07 V_low
+ 1.672010000e-07 V_low
+ 1.673000000e-07 V_low
+ 1.673010000e-07 V_low
+ 1.674000000e-07 V_low
+ 1.674010000e-07 V_low
+ 1.675000000e-07 V_low
+ 1.675010000e-07 V_low
+ 1.676000000e-07 V_low
+ 1.676010000e-07 V_low
+ 1.677000000e-07 V_low
+ 1.677010000e-07 V_low
+ 1.678000000e-07 V_low
+ 1.678010000e-07 V_low
+ 1.679000000e-07 V_low
+ 1.679010000e-07 V_hig
+ 1.680000000e-07 V_hig
+ 1.680010000e-07 V_hig
+ 1.681000000e-07 V_hig
+ 1.681010000e-07 V_hig
+ 1.682000000e-07 V_hig
+ 1.682010000e-07 V_hig
+ 1.683000000e-07 V_hig
+ 1.683010000e-07 V_hig
+ 1.684000000e-07 V_hig
+ 1.684010000e-07 V_hig
+ 1.685000000e-07 V_hig
+ 1.685010000e-07 V_hig
+ 1.686000000e-07 V_hig
+ 1.686010000e-07 V_hig
+ 1.687000000e-07 V_hig
+ 1.687010000e-07 V_hig
+ 1.688000000e-07 V_hig
+ 1.688010000e-07 V_hig
+ 1.689000000e-07 V_hig
+ 1.689010000e-07 V_low
+ 1.690000000e-07 V_low
+ 1.690010000e-07 V_low
+ 1.691000000e-07 V_low
+ 1.691010000e-07 V_low
+ 1.692000000e-07 V_low
+ 1.692010000e-07 V_low
+ 1.693000000e-07 V_low
+ 1.693010000e-07 V_low
+ 1.694000000e-07 V_low
+ 1.694010000e-07 V_low
+ 1.695000000e-07 V_low
+ 1.695010000e-07 V_low
+ 1.696000000e-07 V_low
+ 1.696010000e-07 V_low
+ 1.697000000e-07 V_low
+ 1.697010000e-07 V_low
+ 1.698000000e-07 V_low
+ 1.698010000e-07 V_low
+ 1.699000000e-07 V_low
+ 1.699010000e-07 V_low
+ 1.700000000e-07 V_low
+ 1.700010000e-07 V_low
+ 1.701000000e-07 V_low
+ 1.701010000e-07 V_low
+ 1.702000000e-07 V_low
+ 1.702010000e-07 V_low
+ 1.703000000e-07 V_low
+ 1.703010000e-07 V_low
+ 1.704000000e-07 V_low
+ 1.704010000e-07 V_low
+ 1.705000000e-07 V_low
+ 1.705010000e-07 V_low
+ 1.706000000e-07 V_low
+ 1.706010000e-07 V_low
+ 1.707000000e-07 V_low
+ 1.707010000e-07 V_low
+ 1.708000000e-07 V_low
+ 1.708010000e-07 V_low
+ 1.709000000e-07 V_low
+ 1.709010000e-07 V_hig
+ 1.710000000e-07 V_hig
+ 1.710010000e-07 V_hig
+ 1.711000000e-07 V_hig
+ 1.711010000e-07 V_hig
+ 1.712000000e-07 V_hig
+ 1.712010000e-07 V_hig
+ 1.713000000e-07 V_hig
+ 1.713010000e-07 V_hig
+ 1.714000000e-07 V_hig
+ 1.714010000e-07 V_hig
+ 1.715000000e-07 V_hig
+ 1.715010000e-07 V_hig
+ 1.716000000e-07 V_hig
+ 1.716010000e-07 V_hig
+ 1.717000000e-07 V_hig
+ 1.717010000e-07 V_hig
+ 1.718000000e-07 V_hig
+ 1.718010000e-07 V_hig
+ 1.719000000e-07 V_hig
+ 1.719010000e-07 V_hig
+ 1.720000000e-07 V_hig
+ 1.720010000e-07 V_hig
+ 1.721000000e-07 V_hig
+ 1.721010000e-07 V_hig
+ 1.722000000e-07 V_hig
+ 1.722010000e-07 V_hig
+ 1.723000000e-07 V_hig
+ 1.723010000e-07 V_hig
+ 1.724000000e-07 V_hig
+ 1.724010000e-07 V_hig
+ 1.725000000e-07 V_hig
+ 1.725010000e-07 V_hig
+ 1.726000000e-07 V_hig
+ 1.726010000e-07 V_hig
+ 1.727000000e-07 V_hig
+ 1.727010000e-07 V_hig
+ 1.728000000e-07 V_hig
+ 1.728010000e-07 V_hig
+ 1.729000000e-07 V_hig
+ 1.729010000e-07 V_low
+ 1.730000000e-07 V_low
+ 1.730010000e-07 V_low
+ 1.731000000e-07 V_low
+ 1.731010000e-07 V_low
+ 1.732000000e-07 V_low
+ 1.732010000e-07 V_low
+ 1.733000000e-07 V_low
+ 1.733010000e-07 V_low
+ 1.734000000e-07 V_low
+ 1.734010000e-07 V_low
+ 1.735000000e-07 V_low
+ 1.735010000e-07 V_low
+ 1.736000000e-07 V_low
+ 1.736010000e-07 V_low
+ 1.737000000e-07 V_low
+ 1.737010000e-07 V_low
+ 1.738000000e-07 V_low
+ 1.738010000e-07 V_low
+ 1.739000000e-07 V_low
+ 1.739010000e-07 V_hig
+ 1.740000000e-07 V_hig
+ 1.740010000e-07 V_hig
+ 1.741000000e-07 V_hig
+ 1.741010000e-07 V_hig
+ 1.742000000e-07 V_hig
+ 1.742010000e-07 V_hig
+ 1.743000000e-07 V_hig
+ 1.743010000e-07 V_hig
+ 1.744000000e-07 V_hig
+ 1.744010000e-07 V_hig
+ 1.745000000e-07 V_hig
+ 1.745010000e-07 V_hig
+ 1.746000000e-07 V_hig
+ 1.746010000e-07 V_hig
+ 1.747000000e-07 V_hig
+ 1.747010000e-07 V_hig
+ 1.748000000e-07 V_hig
+ 1.748010000e-07 V_hig
+ 1.749000000e-07 V_hig
+ 1.749010000e-07 V_low
+ 1.750000000e-07 V_low
+ 1.750010000e-07 V_low
+ 1.751000000e-07 V_low
+ 1.751010000e-07 V_low
+ 1.752000000e-07 V_low
+ 1.752010000e-07 V_low
+ 1.753000000e-07 V_low
+ 1.753010000e-07 V_low
+ 1.754000000e-07 V_low
+ 1.754010000e-07 V_low
+ 1.755000000e-07 V_low
+ 1.755010000e-07 V_low
+ 1.756000000e-07 V_low
+ 1.756010000e-07 V_low
+ 1.757000000e-07 V_low
+ 1.757010000e-07 V_low
+ 1.758000000e-07 V_low
+ 1.758010000e-07 V_low
+ 1.759000000e-07 V_low
+ 1.759010000e-07 V_hig
+ 1.760000000e-07 V_hig
+ 1.760010000e-07 V_hig
+ 1.761000000e-07 V_hig
+ 1.761010000e-07 V_hig
+ 1.762000000e-07 V_hig
+ 1.762010000e-07 V_hig
+ 1.763000000e-07 V_hig
+ 1.763010000e-07 V_hig
+ 1.764000000e-07 V_hig
+ 1.764010000e-07 V_hig
+ 1.765000000e-07 V_hig
+ 1.765010000e-07 V_hig
+ 1.766000000e-07 V_hig
+ 1.766010000e-07 V_hig
+ 1.767000000e-07 V_hig
+ 1.767010000e-07 V_hig
+ 1.768000000e-07 V_hig
+ 1.768010000e-07 V_hig
+ 1.769000000e-07 V_hig
+ 1.769010000e-07 V_hig
+ 1.770000000e-07 V_hig
+ 1.770010000e-07 V_hig
+ 1.771000000e-07 V_hig
+ 1.771010000e-07 V_hig
+ 1.772000000e-07 V_hig
+ 1.772010000e-07 V_hig
+ 1.773000000e-07 V_hig
+ 1.773010000e-07 V_hig
+ 1.774000000e-07 V_hig
+ 1.774010000e-07 V_hig
+ 1.775000000e-07 V_hig
+ 1.775010000e-07 V_hig
+ 1.776000000e-07 V_hig
+ 1.776010000e-07 V_hig
+ 1.777000000e-07 V_hig
+ 1.777010000e-07 V_hig
+ 1.778000000e-07 V_hig
+ 1.778010000e-07 V_hig
+ 1.779000000e-07 V_hig
+ 1.779010000e-07 V_hig
+ 1.780000000e-07 V_hig
+ 1.780010000e-07 V_hig
+ 1.781000000e-07 V_hig
+ 1.781010000e-07 V_hig
+ 1.782000000e-07 V_hig
+ 1.782010000e-07 V_hig
+ 1.783000000e-07 V_hig
+ 1.783010000e-07 V_hig
+ 1.784000000e-07 V_hig
+ 1.784010000e-07 V_hig
+ 1.785000000e-07 V_hig
+ 1.785010000e-07 V_hig
+ 1.786000000e-07 V_hig
+ 1.786010000e-07 V_hig
+ 1.787000000e-07 V_hig
+ 1.787010000e-07 V_hig
+ 1.788000000e-07 V_hig
+ 1.788010000e-07 V_hig
+ 1.789000000e-07 V_hig
+ 1.789010000e-07 V_hig
+ 1.790000000e-07 V_hig
+ 1.790010000e-07 V_hig
+ 1.791000000e-07 V_hig
+ 1.791010000e-07 V_hig
+ 1.792000000e-07 V_hig
+ 1.792010000e-07 V_hig
+ 1.793000000e-07 V_hig
+ 1.793010000e-07 V_hig
+ 1.794000000e-07 V_hig
+ 1.794010000e-07 V_hig
+ 1.795000000e-07 V_hig
+ 1.795010000e-07 V_hig
+ 1.796000000e-07 V_hig
+ 1.796010000e-07 V_hig
+ 1.797000000e-07 V_hig
+ 1.797010000e-07 V_hig
+ 1.798000000e-07 V_hig
+ 1.798010000e-07 V_hig
+ 1.799000000e-07 V_hig
+ 1.799010000e-07 V_hig
+ 1.800000000e-07 V_hig
+ 1.800010000e-07 V_hig
+ 1.801000000e-07 V_hig
+ 1.801010000e-07 V_hig
+ 1.802000000e-07 V_hig
+ 1.802010000e-07 V_hig
+ 1.803000000e-07 V_hig
+ 1.803010000e-07 V_hig
+ 1.804000000e-07 V_hig
+ 1.804010000e-07 V_hig
+ 1.805000000e-07 V_hig
+ 1.805010000e-07 V_hig
+ 1.806000000e-07 V_hig
+ 1.806010000e-07 V_hig
+ 1.807000000e-07 V_hig
+ 1.807010000e-07 V_hig
+ 1.808000000e-07 V_hig
+ 1.808010000e-07 V_hig
+ 1.809000000e-07 V_hig
+ 1.809010000e-07 V_hig
+ 1.810000000e-07 V_hig
+ 1.810010000e-07 V_hig
+ 1.811000000e-07 V_hig
+ 1.811010000e-07 V_hig
+ 1.812000000e-07 V_hig
+ 1.812010000e-07 V_hig
+ 1.813000000e-07 V_hig
+ 1.813010000e-07 V_hig
+ 1.814000000e-07 V_hig
+ 1.814010000e-07 V_hig
+ 1.815000000e-07 V_hig
+ 1.815010000e-07 V_hig
+ 1.816000000e-07 V_hig
+ 1.816010000e-07 V_hig
+ 1.817000000e-07 V_hig
+ 1.817010000e-07 V_hig
+ 1.818000000e-07 V_hig
+ 1.818010000e-07 V_hig
+ 1.819000000e-07 V_hig
+ 1.819010000e-07 V_hig
+ 1.820000000e-07 V_hig
+ 1.820010000e-07 V_hig
+ 1.821000000e-07 V_hig
+ 1.821010000e-07 V_hig
+ 1.822000000e-07 V_hig
+ 1.822010000e-07 V_hig
+ 1.823000000e-07 V_hig
+ 1.823010000e-07 V_hig
+ 1.824000000e-07 V_hig
+ 1.824010000e-07 V_hig
+ 1.825000000e-07 V_hig
+ 1.825010000e-07 V_hig
+ 1.826000000e-07 V_hig
+ 1.826010000e-07 V_hig
+ 1.827000000e-07 V_hig
+ 1.827010000e-07 V_hig
+ 1.828000000e-07 V_hig
+ 1.828010000e-07 V_hig
+ 1.829000000e-07 V_hig
+ 1.829010000e-07 V_hig
+ 1.830000000e-07 V_hig
+ 1.830010000e-07 V_hig
+ 1.831000000e-07 V_hig
+ 1.831010000e-07 V_hig
+ 1.832000000e-07 V_hig
+ 1.832010000e-07 V_hig
+ 1.833000000e-07 V_hig
+ 1.833010000e-07 V_hig
+ 1.834000000e-07 V_hig
+ 1.834010000e-07 V_hig
+ 1.835000000e-07 V_hig
+ 1.835010000e-07 V_hig
+ 1.836000000e-07 V_hig
+ 1.836010000e-07 V_hig
+ 1.837000000e-07 V_hig
+ 1.837010000e-07 V_hig
+ 1.838000000e-07 V_hig
+ 1.838010000e-07 V_hig
+ 1.839000000e-07 V_hig
+ 1.839010000e-07 V_hig
+ 1.840000000e-07 V_hig
+ 1.840010000e-07 V_hig
+ 1.841000000e-07 V_hig
+ 1.841010000e-07 V_hig
+ 1.842000000e-07 V_hig
+ 1.842010000e-07 V_hig
+ 1.843000000e-07 V_hig
+ 1.843010000e-07 V_hig
+ 1.844000000e-07 V_hig
+ 1.844010000e-07 V_hig
+ 1.845000000e-07 V_hig
+ 1.845010000e-07 V_hig
+ 1.846000000e-07 V_hig
+ 1.846010000e-07 V_hig
+ 1.847000000e-07 V_hig
+ 1.847010000e-07 V_hig
+ 1.848000000e-07 V_hig
+ 1.848010000e-07 V_hig
+ 1.849000000e-07 V_hig
+ 1.849010000e-07 V_low
+ 1.850000000e-07 V_low
+ 1.850010000e-07 V_low
+ 1.851000000e-07 V_low
+ 1.851010000e-07 V_low
+ 1.852000000e-07 V_low
+ 1.852010000e-07 V_low
+ 1.853000000e-07 V_low
+ 1.853010000e-07 V_low
+ 1.854000000e-07 V_low
+ 1.854010000e-07 V_low
+ 1.855000000e-07 V_low
+ 1.855010000e-07 V_low
+ 1.856000000e-07 V_low
+ 1.856010000e-07 V_low
+ 1.857000000e-07 V_low
+ 1.857010000e-07 V_low
+ 1.858000000e-07 V_low
+ 1.858010000e-07 V_low
+ 1.859000000e-07 V_low
+ 1.859010000e-07 V_hig
+ 1.860000000e-07 V_hig
+ 1.860010000e-07 V_hig
+ 1.861000000e-07 V_hig
+ 1.861010000e-07 V_hig
+ 1.862000000e-07 V_hig
+ 1.862010000e-07 V_hig
+ 1.863000000e-07 V_hig
+ 1.863010000e-07 V_hig
+ 1.864000000e-07 V_hig
+ 1.864010000e-07 V_hig
+ 1.865000000e-07 V_hig
+ 1.865010000e-07 V_hig
+ 1.866000000e-07 V_hig
+ 1.866010000e-07 V_hig
+ 1.867000000e-07 V_hig
+ 1.867010000e-07 V_hig
+ 1.868000000e-07 V_hig
+ 1.868010000e-07 V_hig
+ 1.869000000e-07 V_hig
+ 1.869010000e-07 V_hig
+ 1.870000000e-07 V_hig
+ 1.870010000e-07 V_hig
+ 1.871000000e-07 V_hig
+ 1.871010000e-07 V_hig
+ 1.872000000e-07 V_hig
+ 1.872010000e-07 V_hig
+ 1.873000000e-07 V_hig
+ 1.873010000e-07 V_hig
+ 1.874000000e-07 V_hig
+ 1.874010000e-07 V_hig
+ 1.875000000e-07 V_hig
+ 1.875010000e-07 V_hig
+ 1.876000000e-07 V_hig
+ 1.876010000e-07 V_hig
+ 1.877000000e-07 V_hig
+ 1.877010000e-07 V_hig
+ 1.878000000e-07 V_hig
+ 1.878010000e-07 V_hig
+ 1.879000000e-07 V_hig
+ 1.879010000e-07 V_low
+ 1.880000000e-07 V_low
+ 1.880010000e-07 V_low
+ 1.881000000e-07 V_low
+ 1.881010000e-07 V_low
+ 1.882000000e-07 V_low
+ 1.882010000e-07 V_low
+ 1.883000000e-07 V_low
+ 1.883010000e-07 V_low
+ 1.884000000e-07 V_low
+ 1.884010000e-07 V_low
+ 1.885000000e-07 V_low
+ 1.885010000e-07 V_low
+ 1.886000000e-07 V_low
+ 1.886010000e-07 V_low
+ 1.887000000e-07 V_low
+ 1.887010000e-07 V_low
+ 1.888000000e-07 V_low
+ 1.888010000e-07 V_low
+ 1.889000000e-07 V_low
+ 1.889010000e-07 V_hig
+ 1.890000000e-07 V_hig
+ 1.890010000e-07 V_hig
+ 1.891000000e-07 V_hig
+ 1.891010000e-07 V_hig
+ 1.892000000e-07 V_hig
+ 1.892010000e-07 V_hig
+ 1.893000000e-07 V_hig
+ 1.893010000e-07 V_hig
+ 1.894000000e-07 V_hig
+ 1.894010000e-07 V_hig
+ 1.895000000e-07 V_hig
+ 1.895010000e-07 V_hig
+ 1.896000000e-07 V_hig
+ 1.896010000e-07 V_hig
+ 1.897000000e-07 V_hig
+ 1.897010000e-07 V_hig
+ 1.898000000e-07 V_hig
+ 1.898010000e-07 V_hig
+ 1.899000000e-07 V_hig
+ 1.899010000e-07 V_low
+ 1.900000000e-07 V_low
+ 1.900010000e-07 V_low
+ 1.901000000e-07 V_low
+ 1.901010000e-07 V_low
+ 1.902000000e-07 V_low
+ 1.902010000e-07 V_low
+ 1.903000000e-07 V_low
+ 1.903010000e-07 V_low
+ 1.904000000e-07 V_low
+ 1.904010000e-07 V_low
+ 1.905000000e-07 V_low
+ 1.905010000e-07 V_low
+ 1.906000000e-07 V_low
+ 1.906010000e-07 V_low
+ 1.907000000e-07 V_low
+ 1.907010000e-07 V_low
+ 1.908000000e-07 V_low
+ 1.908010000e-07 V_low
+ 1.909000000e-07 V_low
+ 1.909010000e-07 V_hig
+ 1.910000000e-07 V_hig
+ 1.910010000e-07 V_hig
+ 1.911000000e-07 V_hig
+ 1.911010000e-07 V_hig
+ 1.912000000e-07 V_hig
+ 1.912010000e-07 V_hig
+ 1.913000000e-07 V_hig
+ 1.913010000e-07 V_hig
+ 1.914000000e-07 V_hig
+ 1.914010000e-07 V_hig
+ 1.915000000e-07 V_hig
+ 1.915010000e-07 V_hig
+ 1.916000000e-07 V_hig
+ 1.916010000e-07 V_hig
+ 1.917000000e-07 V_hig
+ 1.917010000e-07 V_hig
+ 1.918000000e-07 V_hig
+ 1.918010000e-07 V_hig
+ 1.919000000e-07 V_hig
+ 1.919010000e-07 V_low
+ 1.920000000e-07 V_low
+ 1.920010000e-07 V_low
+ 1.921000000e-07 V_low
+ 1.921010000e-07 V_low
+ 1.922000000e-07 V_low
+ 1.922010000e-07 V_low
+ 1.923000000e-07 V_low
+ 1.923010000e-07 V_low
+ 1.924000000e-07 V_low
+ 1.924010000e-07 V_low
+ 1.925000000e-07 V_low
+ 1.925010000e-07 V_low
+ 1.926000000e-07 V_low
+ 1.926010000e-07 V_low
+ 1.927000000e-07 V_low
+ 1.927010000e-07 V_low
+ 1.928000000e-07 V_low
+ 1.928010000e-07 V_low
+ 1.929000000e-07 V_low
+ 1.929010000e-07 V_hig
+ 1.930000000e-07 V_hig
+ 1.930010000e-07 V_hig
+ 1.931000000e-07 V_hig
+ 1.931010000e-07 V_hig
+ 1.932000000e-07 V_hig
+ 1.932010000e-07 V_hig
+ 1.933000000e-07 V_hig
+ 1.933010000e-07 V_hig
+ 1.934000000e-07 V_hig
+ 1.934010000e-07 V_hig
+ 1.935000000e-07 V_hig
+ 1.935010000e-07 V_hig
+ 1.936000000e-07 V_hig
+ 1.936010000e-07 V_hig
+ 1.937000000e-07 V_hig
+ 1.937010000e-07 V_hig
+ 1.938000000e-07 V_hig
+ 1.938010000e-07 V_hig
+ 1.939000000e-07 V_hig
+ 1.939010000e-07 V_hig
+ 1.940000000e-07 V_hig
+ 1.940010000e-07 V_hig
+ 1.941000000e-07 V_hig
+ 1.941010000e-07 V_hig
+ 1.942000000e-07 V_hig
+ 1.942010000e-07 V_hig
+ 1.943000000e-07 V_hig
+ 1.943010000e-07 V_hig
+ 1.944000000e-07 V_hig
+ 1.944010000e-07 V_hig
+ 1.945000000e-07 V_hig
+ 1.945010000e-07 V_hig
+ 1.946000000e-07 V_hig
+ 1.946010000e-07 V_hig
+ 1.947000000e-07 V_hig
+ 1.947010000e-07 V_hig
+ 1.948000000e-07 V_hig
+ 1.948010000e-07 V_hig
+ 1.949000000e-07 V_hig
+ 1.949010000e-07 V_low
+ 1.950000000e-07 V_low
+ 1.950010000e-07 V_low
+ 1.951000000e-07 V_low
+ 1.951010000e-07 V_low
+ 1.952000000e-07 V_low
+ 1.952010000e-07 V_low
+ 1.953000000e-07 V_low
+ 1.953010000e-07 V_low
+ 1.954000000e-07 V_low
+ 1.954010000e-07 V_low
+ 1.955000000e-07 V_low
+ 1.955010000e-07 V_low
+ 1.956000000e-07 V_low
+ 1.956010000e-07 V_low
+ 1.957000000e-07 V_low
+ 1.957010000e-07 V_low
+ 1.958000000e-07 V_low
+ 1.958010000e-07 V_low
+ 1.959000000e-07 V_low
+ 1.959010000e-07 V_hig
+ 1.960000000e-07 V_hig
+ 1.960010000e-07 V_hig
+ 1.961000000e-07 V_hig
+ 1.961010000e-07 V_hig
+ 1.962000000e-07 V_hig
+ 1.962010000e-07 V_hig
+ 1.963000000e-07 V_hig
+ 1.963010000e-07 V_hig
+ 1.964000000e-07 V_hig
+ 1.964010000e-07 V_hig
+ 1.965000000e-07 V_hig
+ 1.965010000e-07 V_hig
+ 1.966000000e-07 V_hig
+ 1.966010000e-07 V_hig
+ 1.967000000e-07 V_hig
+ 1.967010000e-07 V_hig
+ 1.968000000e-07 V_hig
+ 1.968010000e-07 V_hig
+ 1.969000000e-07 V_hig
+ 1.969010000e-07 V_hig
+ 1.970000000e-07 V_hig
+ 1.970010000e-07 V_hig
+ 1.971000000e-07 V_hig
+ 1.971010000e-07 V_hig
+ 1.972000000e-07 V_hig
+ 1.972010000e-07 V_hig
+ 1.973000000e-07 V_hig
+ 1.973010000e-07 V_hig
+ 1.974000000e-07 V_hig
+ 1.974010000e-07 V_hig
+ 1.975000000e-07 V_hig
+ 1.975010000e-07 V_hig
+ 1.976000000e-07 V_hig
+ 1.976010000e-07 V_hig
+ 1.977000000e-07 V_hig
+ 1.977010000e-07 V_hig
+ 1.978000000e-07 V_hig
+ 1.978010000e-07 V_hig
+ 1.979000000e-07 V_hig
+ 1.979010000e-07 V_low
+ 1.980000000e-07 V_low
+ 1.980010000e-07 V_low
+ 1.981000000e-07 V_low
+ 1.981010000e-07 V_low
+ 1.982000000e-07 V_low
+ 1.982010000e-07 V_low
+ 1.983000000e-07 V_low
+ 1.983010000e-07 V_low
+ 1.984000000e-07 V_low
+ 1.984010000e-07 V_low
+ 1.985000000e-07 V_low
+ 1.985010000e-07 V_low
+ 1.986000000e-07 V_low
+ 1.986010000e-07 V_low
+ 1.987000000e-07 V_low
+ 1.987010000e-07 V_low
+ 1.988000000e-07 V_low
+ 1.988010000e-07 V_low
+ 1.989000000e-07 V_low
+ 1.989010000e-07 V_hig
+ 1.990000000e-07 V_hig
+ 1.990010000e-07 V_hig
+ 1.991000000e-07 V_hig
+ 1.991010000e-07 V_hig
+ 1.992000000e-07 V_hig
+ 1.992010000e-07 V_hig
+ 1.993000000e-07 V_hig
+ 1.993010000e-07 V_hig
+ 1.994000000e-07 V_hig
+ 1.994010000e-07 V_hig
+ 1.995000000e-07 V_hig
+ 1.995010000e-07 V_hig
+ 1.996000000e-07 V_hig
+ 1.996010000e-07 V_hig
+ 1.997000000e-07 V_hig
+ 1.997010000e-07 V_hig
+ 1.998000000e-07 V_hig
+ 1.998010000e-07 V_hig
+ 1.999000000e-07 V_hig
+ 1.999010000e-07 V_hig
+ 2.000000000e-07 V_hig
+ 2.000010000e-07 V_hig
+ 2.001000000e-07 V_hig
+ 2.001010000e-07 V_hig
+ 2.002000000e-07 V_hig
+ 2.002010000e-07 V_hig
+ 2.003000000e-07 V_hig
+ 2.003010000e-07 V_hig
+ 2.004000000e-07 V_hig
+ 2.004010000e-07 V_hig
+ 2.005000000e-07 V_hig
+ 2.005010000e-07 V_hig
+ 2.006000000e-07 V_hig
+ 2.006010000e-07 V_hig
+ 2.007000000e-07 V_hig
+ 2.007010000e-07 V_hig
+ 2.008000000e-07 V_hig
+ 2.008010000e-07 V_hig
+ 2.009000000e-07 V_hig
+ 2.009010000e-07 V_low
+ 2.010000000e-07 V_low
+ 2.010010000e-07 V_low
+ 2.011000000e-07 V_low
+ 2.011010000e-07 V_low
+ 2.012000000e-07 V_low
+ 2.012010000e-07 V_low
+ 2.013000000e-07 V_low
+ 2.013010000e-07 V_low
+ 2.014000000e-07 V_low
+ 2.014010000e-07 V_low
+ 2.015000000e-07 V_low
+ 2.015010000e-07 V_low
+ 2.016000000e-07 V_low
+ 2.016010000e-07 V_low
+ 2.017000000e-07 V_low
+ 2.017010000e-07 V_low
+ 2.018000000e-07 V_low
+ 2.018010000e-07 V_low
+ 2.019000000e-07 V_low
+ 2.019010000e-07 V_hig
+ 2.020000000e-07 V_hig
+ 2.020010000e-07 V_hig
+ 2.021000000e-07 V_hig
+ 2.021010000e-07 V_hig
+ 2.022000000e-07 V_hig
+ 2.022010000e-07 V_hig
+ 2.023000000e-07 V_hig
+ 2.023010000e-07 V_hig
+ 2.024000000e-07 V_hig
+ 2.024010000e-07 V_hig
+ 2.025000000e-07 V_hig
+ 2.025010000e-07 V_hig
+ 2.026000000e-07 V_hig
+ 2.026010000e-07 V_hig
+ 2.027000000e-07 V_hig
+ 2.027010000e-07 V_hig
+ 2.028000000e-07 V_hig
+ 2.028010000e-07 V_hig
+ 2.029000000e-07 V_hig
+ 2.029010000e-07 V_hig
+ 2.030000000e-07 V_hig
+ 2.030010000e-07 V_hig
+ 2.031000000e-07 V_hig
+ 2.031010000e-07 V_hig
+ 2.032000000e-07 V_hig
+ 2.032010000e-07 V_hig
+ 2.033000000e-07 V_hig
+ 2.033010000e-07 V_hig
+ 2.034000000e-07 V_hig
+ 2.034010000e-07 V_hig
+ 2.035000000e-07 V_hig
+ 2.035010000e-07 V_hig
+ 2.036000000e-07 V_hig
+ 2.036010000e-07 V_hig
+ 2.037000000e-07 V_hig
+ 2.037010000e-07 V_hig
+ 2.038000000e-07 V_hig
+ 2.038010000e-07 V_hig
+ 2.039000000e-07 V_hig
+ 2.039010000e-07 V_hig
+ 2.040000000e-07 V_hig
+ 2.040010000e-07 V_hig
+ 2.041000000e-07 V_hig
+ 2.041010000e-07 V_hig
+ 2.042000000e-07 V_hig
+ 2.042010000e-07 V_hig
+ 2.043000000e-07 V_hig
+ 2.043010000e-07 V_hig
+ 2.044000000e-07 V_hig
+ 2.044010000e-07 V_hig
+ 2.045000000e-07 V_hig
+ 2.045010000e-07 V_hig
+ 2.046000000e-07 V_hig
+ 2.046010000e-07 V_hig
+ 2.047000000e-07 V_hig
+ 2.047010000e-07 V_hig
+ 2.048000000e-07 V_hig
+ 2.048010000e-07 V_hig
+ 2.049000000e-07 V_hig
+ 2.049010000e-07 V_hig
+ 2.050000000e-07 V_hig
+ 2.050010000e-07 V_hig
+ 2.051000000e-07 V_hig
+ 2.051010000e-07 V_hig
+ 2.052000000e-07 V_hig
+ 2.052010000e-07 V_hig
+ 2.053000000e-07 V_hig
+ 2.053010000e-07 V_hig
+ 2.054000000e-07 V_hig
+ 2.054010000e-07 V_hig
+ 2.055000000e-07 V_hig
+ 2.055010000e-07 V_hig
+ 2.056000000e-07 V_hig
+ 2.056010000e-07 V_hig
+ 2.057000000e-07 V_hig
+ 2.057010000e-07 V_hig
+ 2.058000000e-07 V_hig
+ 2.058010000e-07 V_hig
+ 2.059000000e-07 V_hig
+ 2.059010000e-07 V_low
+ 2.060000000e-07 V_low
+ 2.060010000e-07 V_low
+ 2.061000000e-07 V_low
+ 2.061010000e-07 V_low
+ 2.062000000e-07 V_low
+ 2.062010000e-07 V_low
+ 2.063000000e-07 V_low
+ 2.063010000e-07 V_low
+ 2.064000000e-07 V_low
+ 2.064010000e-07 V_low
+ 2.065000000e-07 V_low
+ 2.065010000e-07 V_low
+ 2.066000000e-07 V_low
+ 2.066010000e-07 V_low
+ 2.067000000e-07 V_low
+ 2.067010000e-07 V_low
+ 2.068000000e-07 V_low
+ 2.068010000e-07 V_low
+ 2.069000000e-07 V_low
+ 2.069010000e-07 V_low
+ 2.070000000e-07 V_low
+ 2.070010000e-07 V_low
+ 2.071000000e-07 V_low
+ 2.071010000e-07 V_low
+ 2.072000000e-07 V_low
+ 2.072010000e-07 V_low
+ 2.073000000e-07 V_low
+ 2.073010000e-07 V_low
+ 2.074000000e-07 V_low
+ 2.074010000e-07 V_low
+ 2.075000000e-07 V_low
+ 2.075010000e-07 V_low
+ 2.076000000e-07 V_low
+ 2.076010000e-07 V_low
+ 2.077000000e-07 V_low
+ 2.077010000e-07 V_low
+ 2.078000000e-07 V_low
+ 2.078010000e-07 V_low
+ 2.079000000e-07 V_low
+ 2.079010000e-07 V_hig
+ 2.080000000e-07 V_hig
+ 2.080010000e-07 V_hig
+ 2.081000000e-07 V_hig
+ 2.081010000e-07 V_hig
+ 2.082000000e-07 V_hig
+ 2.082010000e-07 V_hig
+ 2.083000000e-07 V_hig
+ 2.083010000e-07 V_hig
+ 2.084000000e-07 V_hig
+ 2.084010000e-07 V_hig
+ 2.085000000e-07 V_hig
+ 2.085010000e-07 V_hig
+ 2.086000000e-07 V_hig
+ 2.086010000e-07 V_hig
+ 2.087000000e-07 V_hig
+ 2.087010000e-07 V_hig
+ 2.088000000e-07 V_hig
+ 2.088010000e-07 V_hig
+ 2.089000000e-07 V_hig
+ 2.089010000e-07 V_low
+ 2.090000000e-07 V_low
+ 2.090010000e-07 V_low
+ 2.091000000e-07 V_low
+ 2.091010000e-07 V_low
+ 2.092000000e-07 V_low
+ 2.092010000e-07 V_low
+ 2.093000000e-07 V_low
+ 2.093010000e-07 V_low
+ 2.094000000e-07 V_low
+ 2.094010000e-07 V_low
+ 2.095000000e-07 V_low
+ 2.095010000e-07 V_low
+ 2.096000000e-07 V_low
+ 2.096010000e-07 V_low
+ 2.097000000e-07 V_low
+ 2.097010000e-07 V_low
+ 2.098000000e-07 V_low
+ 2.098010000e-07 V_low
+ 2.099000000e-07 V_low
+ 2.099010000e-07 V_low
+ 2.100000000e-07 V_low
+ 2.100010000e-07 V_low
+ 2.101000000e-07 V_low
+ 2.101010000e-07 V_low
+ 2.102000000e-07 V_low
+ 2.102010000e-07 V_low
+ 2.103000000e-07 V_low
+ 2.103010000e-07 V_low
+ 2.104000000e-07 V_low
+ 2.104010000e-07 V_low
+ 2.105000000e-07 V_low
+ 2.105010000e-07 V_low
+ 2.106000000e-07 V_low
+ 2.106010000e-07 V_low
+ 2.107000000e-07 V_low
+ 2.107010000e-07 V_low
+ 2.108000000e-07 V_low
+ 2.108010000e-07 V_low
+ 2.109000000e-07 V_low
+ 2.109010000e-07 V_hig
+ 2.110000000e-07 V_hig
+ 2.110010000e-07 V_hig
+ 2.111000000e-07 V_hig
+ 2.111010000e-07 V_hig
+ 2.112000000e-07 V_hig
+ 2.112010000e-07 V_hig
+ 2.113000000e-07 V_hig
+ 2.113010000e-07 V_hig
+ 2.114000000e-07 V_hig
+ 2.114010000e-07 V_hig
+ 2.115000000e-07 V_hig
+ 2.115010000e-07 V_hig
+ 2.116000000e-07 V_hig
+ 2.116010000e-07 V_hig
+ 2.117000000e-07 V_hig
+ 2.117010000e-07 V_hig
+ 2.118000000e-07 V_hig
+ 2.118010000e-07 V_hig
+ 2.119000000e-07 V_hig
+ 2.119010000e-07 V_low
+ 2.120000000e-07 V_low
+ 2.120010000e-07 V_low
+ 2.121000000e-07 V_low
+ 2.121010000e-07 V_low
+ 2.122000000e-07 V_low
+ 2.122010000e-07 V_low
+ 2.123000000e-07 V_low
+ 2.123010000e-07 V_low
+ 2.124000000e-07 V_low
+ 2.124010000e-07 V_low
+ 2.125000000e-07 V_low
+ 2.125010000e-07 V_low
+ 2.126000000e-07 V_low
+ 2.126010000e-07 V_low
+ 2.127000000e-07 V_low
+ 2.127010000e-07 V_low
+ 2.128000000e-07 V_low
+ 2.128010000e-07 V_low
+ 2.129000000e-07 V_low
+ 2.129010000e-07 V_low
+ 2.130000000e-07 V_low
+ 2.130010000e-07 V_low
+ 2.131000000e-07 V_low
+ 2.131010000e-07 V_low
+ 2.132000000e-07 V_low
+ 2.132010000e-07 V_low
+ 2.133000000e-07 V_low
+ 2.133010000e-07 V_low
+ 2.134000000e-07 V_low
+ 2.134010000e-07 V_low
+ 2.135000000e-07 V_low
+ 2.135010000e-07 V_low
+ 2.136000000e-07 V_low
+ 2.136010000e-07 V_low
+ 2.137000000e-07 V_low
+ 2.137010000e-07 V_low
+ 2.138000000e-07 V_low
+ 2.138010000e-07 V_low
+ 2.139000000e-07 V_low
+ 2.139010000e-07 V_hig
+ 2.140000000e-07 V_hig
+ 2.140010000e-07 V_hig
+ 2.141000000e-07 V_hig
+ 2.141010000e-07 V_hig
+ 2.142000000e-07 V_hig
+ 2.142010000e-07 V_hig
+ 2.143000000e-07 V_hig
+ 2.143010000e-07 V_hig
+ 2.144000000e-07 V_hig
+ 2.144010000e-07 V_hig
+ 2.145000000e-07 V_hig
+ 2.145010000e-07 V_hig
+ 2.146000000e-07 V_hig
+ 2.146010000e-07 V_hig
+ 2.147000000e-07 V_hig
+ 2.147010000e-07 V_hig
+ 2.148000000e-07 V_hig
+ 2.148010000e-07 V_hig
+ 2.149000000e-07 V_hig
+ 2.149010000e-07 V_low
+ 2.150000000e-07 V_low
+ 2.150010000e-07 V_low
+ 2.151000000e-07 V_low
+ 2.151010000e-07 V_low
+ 2.152000000e-07 V_low
+ 2.152010000e-07 V_low
+ 2.153000000e-07 V_low
+ 2.153010000e-07 V_low
+ 2.154000000e-07 V_low
+ 2.154010000e-07 V_low
+ 2.155000000e-07 V_low
+ 2.155010000e-07 V_low
+ 2.156000000e-07 V_low
+ 2.156010000e-07 V_low
+ 2.157000000e-07 V_low
+ 2.157010000e-07 V_low
+ 2.158000000e-07 V_low
+ 2.158010000e-07 V_low
+ 2.159000000e-07 V_low
+ 2.159010000e-07 V_hig
+ 2.160000000e-07 V_hig
+ 2.160010000e-07 V_hig
+ 2.161000000e-07 V_hig
+ 2.161010000e-07 V_hig
+ 2.162000000e-07 V_hig
+ 2.162010000e-07 V_hig
+ 2.163000000e-07 V_hig
+ 2.163010000e-07 V_hig
+ 2.164000000e-07 V_hig
+ 2.164010000e-07 V_hig
+ 2.165000000e-07 V_hig
+ 2.165010000e-07 V_hig
+ 2.166000000e-07 V_hig
+ 2.166010000e-07 V_hig
+ 2.167000000e-07 V_hig
+ 2.167010000e-07 V_hig
+ 2.168000000e-07 V_hig
+ 2.168010000e-07 V_hig
+ 2.169000000e-07 V_hig
+ 2.169010000e-07 V_low
+ 2.170000000e-07 V_low
+ 2.170010000e-07 V_low
+ 2.171000000e-07 V_low
+ 2.171010000e-07 V_low
+ 2.172000000e-07 V_low
+ 2.172010000e-07 V_low
+ 2.173000000e-07 V_low
+ 2.173010000e-07 V_low
+ 2.174000000e-07 V_low
+ 2.174010000e-07 V_low
+ 2.175000000e-07 V_low
+ 2.175010000e-07 V_low
+ 2.176000000e-07 V_low
+ 2.176010000e-07 V_low
+ 2.177000000e-07 V_low
+ 2.177010000e-07 V_low
+ 2.178000000e-07 V_low
+ 2.178010000e-07 V_low
+ 2.179000000e-07 V_low
+ 2.179010000e-07 V_low
+ 2.180000000e-07 V_low
+ 2.180010000e-07 V_low
+ 2.181000000e-07 V_low
+ 2.181010000e-07 V_low
+ 2.182000000e-07 V_low
+ 2.182010000e-07 V_low
+ 2.183000000e-07 V_low
+ 2.183010000e-07 V_low
+ 2.184000000e-07 V_low
+ 2.184010000e-07 V_low
+ 2.185000000e-07 V_low
+ 2.185010000e-07 V_low
+ 2.186000000e-07 V_low
+ 2.186010000e-07 V_low
+ 2.187000000e-07 V_low
+ 2.187010000e-07 V_low
+ 2.188000000e-07 V_low
+ 2.188010000e-07 V_low
+ 2.189000000e-07 V_low
+ 2.189010000e-07 V_low
+ 2.190000000e-07 V_low
+ 2.190010000e-07 V_low
+ 2.191000000e-07 V_low
+ 2.191010000e-07 V_low
+ 2.192000000e-07 V_low
+ 2.192010000e-07 V_low
+ 2.193000000e-07 V_low
+ 2.193010000e-07 V_low
+ 2.194000000e-07 V_low
+ 2.194010000e-07 V_low
+ 2.195000000e-07 V_low
+ 2.195010000e-07 V_low
+ 2.196000000e-07 V_low
+ 2.196010000e-07 V_low
+ 2.197000000e-07 V_low
+ 2.197010000e-07 V_low
+ 2.198000000e-07 V_low
+ 2.198010000e-07 V_low
+ 2.199000000e-07 V_low
+ 2.199010000e-07 V_low
+ 2.200000000e-07 V_low
+ 2.200010000e-07 V_low
+ 2.201000000e-07 V_low
+ 2.201010000e-07 V_low
+ 2.202000000e-07 V_low
+ 2.202010000e-07 V_low
+ 2.203000000e-07 V_low
+ 2.203010000e-07 V_low
+ 2.204000000e-07 V_low
+ 2.204010000e-07 V_low
+ 2.205000000e-07 V_low
+ 2.205010000e-07 V_low
+ 2.206000000e-07 V_low
+ 2.206010000e-07 V_low
+ 2.207000000e-07 V_low
+ 2.207010000e-07 V_low
+ 2.208000000e-07 V_low
+ 2.208010000e-07 V_low
+ 2.209000000e-07 V_low
+ 2.209010000e-07 V_low
+ 2.210000000e-07 V_low
+ 2.210010000e-07 V_low
+ 2.211000000e-07 V_low
+ 2.211010000e-07 V_low
+ 2.212000000e-07 V_low
+ 2.212010000e-07 V_low
+ 2.213000000e-07 V_low
+ 2.213010000e-07 V_low
+ 2.214000000e-07 V_low
+ 2.214010000e-07 V_low
+ 2.215000000e-07 V_low
+ 2.215010000e-07 V_low
+ 2.216000000e-07 V_low
+ 2.216010000e-07 V_low
+ 2.217000000e-07 V_low
+ 2.217010000e-07 V_low
+ 2.218000000e-07 V_low
+ 2.218010000e-07 V_low
+ 2.219000000e-07 V_low
+ 2.219010000e-07 V_hig
+ 2.220000000e-07 V_hig
+ 2.220010000e-07 V_hig
+ 2.221000000e-07 V_hig
+ 2.221010000e-07 V_hig
+ 2.222000000e-07 V_hig
+ 2.222010000e-07 V_hig
+ 2.223000000e-07 V_hig
+ 2.223010000e-07 V_hig
+ 2.224000000e-07 V_hig
+ 2.224010000e-07 V_hig
+ 2.225000000e-07 V_hig
+ 2.225010000e-07 V_hig
+ 2.226000000e-07 V_hig
+ 2.226010000e-07 V_hig
+ 2.227000000e-07 V_hig
+ 2.227010000e-07 V_hig
+ 2.228000000e-07 V_hig
+ 2.228010000e-07 V_hig
+ 2.229000000e-07 V_hig
+ 2.229010000e-07 V_hig
+ 2.230000000e-07 V_hig
+ 2.230010000e-07 V_hig
+ 2.231000000e-07 V_hig
+ 2.231010000e-07 V_hig
+ 2.232000000e-07 V_hig
+ 2.232010000e-07 V_hig
+ 2.233000000e-07 V_hig
+ 2.233010000e-07 V_hig
+ 2.234000000e-07 V_hig
+ 2.234010000e-07 V_hig
+ 2.235000000e-07 V_hig
+ 2.235010000e-07 V_hig
+ 2.236000000e-07 V_hig
+ 2.236010000e-07 V_hig
+ 2.237000000e-07 V_hig
+ 2.237010000e-07 V_hig
+ 2.238000000e-07 V_hig
+ 2.238010000e-07 V_hig
+ 2.239000000e-07 V_hig
+ 2.239010000e-07 V_hig
+ 2.240000000e-07 V_hig
+ 2.240010000e-07 V_hig
+ 2.241000000e-07 V_hig
+ 2.241010000e-07 V_hig
+ 2.242000000e-07 V_hig
+ 2.242010000e-07 V_hig
+ 2.243000000e-07 V_hig
+ 2.243010000e-07 V_hig
+ 2.244000000e-07 V_hig
+ 2.244010000e-07 V_hig
+ 2.245000000e-07 V_hig
+ 2.245010000e-07 V_hig
+ 2.246000000e-07 V_hig
+ 2.246010000e-07 V_hig
+ 2.247000000e-07 V_hig
+ 2.247010000e-07 V_hig
+ 2.248000000e-07 V_hig
+ 2.248010000e-07 V_hig
+ 2.249000000e-07 V_hig
+ 2.249010000e-07 V_hig
+ 2.250000000e-07 V_hig
+ 2.250010000e-07 V_hig
+ 2.251000000e-07 V_hig
+ 2.251010000e-07 V_hig
+ 2.252000000e-07 V_hig
+ 2.252010000e-07 V_hig
+ 2.253000000e-07 V_hig
+ 2.253010000e-07 V_hig
+ 2.254000000e-07 V_hig
+ 2.254010000e-07 V_hig
+ 2.255000000e-07 V_hig
+ 2.255010000e-07 V_hig
+ 2.256000000e-07 V_hig
+ 2.256010000e-07 V_hig
+ 2.257000000e-07 V_hig
+ 2.257010000e-07 V_hig
+ 2.258000000e-07 V_hig
+ 2.258010000e-07 V_hig
+ 2.259000000e-07 V_hig
+ 2.259010000e-07 V_low
+ 2.260000000e-07 V_low
+ 2.260010000e-07 V_low
+ 2.261000000e-07 V_low
+ 2.261010000e-07 V_low
+ 2.262000000e-07 V_low
+ 2.262010000e-07 V_low
+ 2.263000000e-07 V_low
+ 2.263010000e-07 V_low
+ 2.264000000e-07 V_low
+ 2.264010000e-07 V_low
+ 2.265000000e-07 V_low
+ 2.265010000e-07 V_low
+ 2.266000000e-07 V_low
+ 2.266010000e-07 V_low
+ 2.267000000e-07 V_low
+ 2.267010000e-07 V_low
+ 2.268000000e-07 V_low
+ 2.268010000e-07 V_low
+ 2.269000000e-07 V_low
+ 2.269010000e-07 V_low
+ 2.270000000e-07 V_low
+ 2.270010000e-07 V_low
+ 2.271000000e-07 V_low
+ 2.271010000e-07 V_low
+ 2.272000000e-07 V_low
+ 2.272010000e-07 V_low
+ 2.273000000e-07 V_low
+ 2.273010000e-07 V_low
+ 2.274000000e-07 V_low
+ 2.274010000e-07 V_low
+ 2.275000000e-07 V_low
+ 2.275010000e-07 V_low
+ 2.276000000e-07 V_low
+ 2.276010000e-07 V_low
+ 2.277000000e-07 V_low
+ 2.277010000e-07 V_low
+ 2.278000000e-07 V_low
+ 2.278010000e-07 V_low
+ 2.279000000e-07 V_low
+ 2.279010000e-07 V_low
+ 2.280000000e-07 V_low
+ 2.280010000e-07 V_low
+ 2.281000000e-07 V_low
+ 2.281010000e-07 V_low
+ 2.282000000e-07 V_low
+ 2.282010000e-07 V_low
+ 2.283000000e-07 V_low
+ 2.283010000e-07 V_low
+ 2.284000000e-07 V_low
+ 2.284010000e-07 V_low
+ 2.285000000e-07 V_low
+ 2.285010000e-07 V_low
+ 2.286000000e-07 V_low
+ 2.286010000e-07 V_low
+ 2.287000000e-07 V_low
+ 2.287010000e-07 V_low
+ 2.288000000e-07 V_low
+ 2.288010000e-07 V_low
+ 2.289000000e-07 V_low
+ 2.289010000e-07 V_hig
+ 2.290000000e-07 V_hig
+ 2.290010000e-07 V_hig
+ 2.291000000e-07 V_hig
+ 2.291010000e-07 V_hig
+ 2.292000000e-07 V_hig
+ 2.292010000e-07 V_hig
+ 2.293000000e-07 V_hig
+ 2.293010000e-07 V_hig
+ 2.294000000e-07 V_hig
+ 2.294010000e-07 V_hig
+ 2.295000000e-07 V_hig
+ 2.295010000e-07 V_hig
+ 2.296000000e-07 V_hig
+ 2.296010000e-07 V_hig
+ 2.297000000e-07 V_hig
+ 2.297010000e-07 V_hig
+ 2.298000000e-07 V_hig
+ 2.298010000e-07 V_hig
+ 2.299000000e-07 V_hig
+ 2.299010000e-07 V_hig
+ 2.300000000e-07 V_hig
+ 2.300010000e-07 V_hig
+ 2.301000000e-07 V_hig
+ 2.301010000e-07 V_hig
+ 2.302000000e-07 V_hig
+ 2.302010000e-07 V_hig
+ 2.303000000e-07 V_hig
+ 2.303010000e-07 V_hig
+ 2.304000000e-07 V_hig
+ 2.304010000e-07 V_hig
+ 2.305000000e-07 V_hig
+ 2.305010000e-07 V_hig
+ 2.306000000e-07 V_hig
+ 2.306010000e-07 V_hig
+ 2.307000000e-07 V_hig
+ 2.307010000e-07 V_hig
+ 2.308000000e-07 V_hig
+ 2.308010000e-07 V_hig
+ 2.309000000e-07 V_hig
+ 2.309010000e-07 V_hig
+ 2.310000000e-07 V_hig
+ 2.310010000e-07 V_hig
+ 2.311000000e-07 V_hig
+ 2.311010000e-07 V_hig
+ 2.312000000e-07 V_hig
+ 2.312010000e-07 V_hig
+ 2.313000000e-07 V_hig
+ 2.313010000e-07 V_hig
+ 2.314000000e-07 V_hig
+ 2.314010000e-07 V_hig
+ 2.315000000e-07 V_hig
+ 2.315010000e-07 V_hig
+ 2.316000000e-07 V_hig
+ 2.316010000e-07 V_hig
+ 2.317000000e-07 V_hig
+ 2.317010000e-07 V_hig
+ 2.318000000e-07 V_hig
+ 2.318010000e-07 V_hig
+ 2.319000000e-07 V_hig
+ 2.319010000e-07 V_low
+ 2.320000000e-07 V_low
+ 2.320010000e-07 V_low
+ 2.321000000e-07 V_low
+ 2.321010000e-07 V_low
+ 2.322000000e-07 V_low
+ 2.322010000e-07 V_low
+ 2.323000000e-07 V_low
+ 2.323010000e-07 V_low
+ 2.324000000e-07 V_low
+ 2.324010000e-07 V_low
+ 2.325000000e-07 V_low
+ 2.325010000e-07 V_low
+ 2.326000000e-07 V_low
+ 2.326010000e-07 V_low
+ 2.327000000e-07 V_low
+ 2.327010000e-07 V_low
+ 2.328000000e-07 V_low
+ 2.328010000e-07 V_low
+ 2.329000000e-07 V_low
+ 2.329010000e-07 V_hig
+ 2.330000000e-07 V_hig
+ 2.330010000e-07 V_hig
+ 2.331000000e-07 V_hig
+ 2.331010000e-07 V_hig
+ 2.332000000e-07 V_hig
+ 2.332010000e-07 V_hig
+ 2.333000000e-07 V_hig
+ 2.333010000e-07 V_hig
+ 2.334000000e-07 V_hig
+ 2.334010000e-07 V_hig
+ 2.335000000e-07 V_hig
+ 2.335010000e-07 V_hig
+ 2.336000000e-07 V_hig
+ 2.336010000e-07 V_hig
+ 2.337000000e-07 V_hig
+ 2.337010000e-07 V_hig
+ 2.338000000e-07 V_hig
+ 2.338010000e-07 V_hig
+ 2.339000000e-07 V_hig
+ 2.339010000e-07 V_hig
+ 2.340000000e-07 V_hig
+ 2.340010000e-07 V_hig
+ 2.341000000e-07 V_hig
+ 2.341010000e-07 V_hig
+ 2.342000000e-07 V_hig
+ 2.342010000e-07 V_hig
+ 2.343000000e-07 V_hig
+ 2.343010000e-07 V_hig
+ 2.344000000e-07 V_hig
+ 2.344010000e-07 V_hig
+ 2.345000000e-07 V_hig
+ 2.345010000e-07 V_hig
+ 2.346000000e-07 V_hig
+ 2.346010000e-07 V_hig
+ 2.347000000e-07 V_hig
+ 2.347010000e-07 V_hig
+ 2.348000000e-07 V_hig
+ 2.348010000e-07 V_hig
+ 2.349000000e-07 V_hig
+ 2.349010000e-07 V_hig
+ 2.350000000e-07 V_hig
+ 2.350010000e-07 V_hig
+ 2.351000000e-07 V_hig
+ 2.351010000e-07 V_hig
+ 2.352000000e-07 V_hig
+ 2.352010000e-07 V_hig
+ 2.353000000e-07 V_hig
+ 2.353010000e-07 V_hig
+ 2.354000000e-07 V_hig
+ 2.354010000e-07 V_hig
+ 2.355000000e-07 V_hig
+ 2.355010000e-07 V_hig
+ 2.356000000e-07 V_hig
+ 2.356010000e-07 V_hig
+ 2.357000000e-07 V_hig
+ 2.357010000e-07 V_hig
+ 2.358000000e-07 V_hig
+ 2.358010000e-07 V_hig
+ 2.359000000e-07 V_hig
+ 2.359010000e-07 V_hig
+ 2.360000000e-07 V_hig
+ 2.360010000e-07 V_hig
+ 2.361000000e-07 V_hig
+ 2.361010000e-07 V_hig
+ 2.362000000e-07 V_hig
+ 2.362010000e-07 V_hig
+ 2.363000000e-07 V_hig
+ 2.363010000e-07 V_hig
+ 2.364000000e-07 V_hig
+ 2.364010000e-07 V_hig
+ 2.365000000e-07 V_hig
+ 2.365010000e-07 V_hig
+ 2.366000000e-07 V_hig
+ 2.366010000e-07 V_hig
+ 2.367000000e-07 V_hig
+ 2.367010000e-07 V_hig
+ 2.368000000e-07 V_hig
+ 2.368010000e-07 V_hig
+ 2.369000000e-07 V_hig
+ 2.369010000e-07 V_low
+ 2.370000000e-07 V_low
+ 2.370010000e-07 V_low
+ 2.371000000e-07 V_low
+ 2.371010000e-07 V_low
+ 2.372000000e-07 V_low
+ 2.372010000e-07 V_low
+ 2.373000000e-07 V_low
+ 2.373010000e-07 V_low
+ 2.374000000e-07 V_low
+ 2.374010000e-07 V_low
+ 2.375000000e-07 V_low
+ 2.375010000e-07 V_low
+ 2.376000000e-07 V_low
+ 2.376010000e-07 V_low
+ 2.377000000e-07 V_low
+ 2.377010000e-07 V_low
+ 2.378000000e-07 V_low
+ 2.378010000e-07 V_low
+ 2.379000000e-07 V_low
+ 2.379010000e-07 V_hig
+ 2.380000000e-07 V_hig
+ 2.380010000e-07 V_hig
+ 2.381000000e-07 V_hig
+ 2.381010000e-07 V_hig
+ 2.382000000e-07 V_hig
+ 2.382010000e-07 V_hig
+ 2.383000000e-07 V_hig
+ 2.383010000e-07 V_hig
+ 2.384000000e-07 V_hig
+ 2.384010000e-07 V_hig
+ 2.385000000e-07 V_hig
+ 2.385010000e-07 V_hig
+ 2.386000000e-07 V_hig
+ 2.386010000e-07 V_hig
+ 2.387000000e-07 V_hig
+ 2.387010000e-07 V_hig
+ 2.388000000e-07 V_hig
+ 2.388010000e-07 V_hig
+ 2.389000000e-07 V_hig
+ 2.389010000e-07 V_low
+ 2.390000000e-07 V_low
+ 2.390010000e-07 V_low
+ 2.391000000e-07 V_low
+ 2.391010000e-07 V_low
+ 2.392000000e-07 V_low
+ 2.392010000e-07 V_low
+ 2.393000000e-07 V_low
+ 2.393010000e-07 V_low
+ 2.394000000e-07 V_low
+ 2.394010000e-07 V_low
+ 2.395000000e-07 V_low
+ 2.395010000e-07 V_low
+ 2.396000000e-07 V_low
+ 2.396010000e-07 V_low
+ 2.397000000e-07 V_low
+ 2.397010000e-07 V_low
+ 2.398000000e-07 V_low
+ 2.398010000e-07 V_low
+ 2.399000000e-07 V_low
+ 2.399010000e-07 V_hig
+ 2.400000000e-07 V_hig
+ 2.400010000e-07 V_hig
+ 2.401000000e-07 V_hig
+ 2.401010000e-07 V_hig
+ 2.402000000e-07 V_hig
+ 2.402010000e-07 V_hig
+ 2.403000000e-07 V_hig
+ 2.403010000e-07 V_hig
+ 2.404000000e-07 V_hig
+ 2.404010000e-07 V_hig
+ 2.405000000e-07 V_hig
+ 2.405010000e-07 V_hig
+ 2.406000000e-07 V_hig
+ 2.406010000e-07 V_hig
+ 2.407000000e-07 V_hig
+ 2.407010000e-07 V_hig
+ 2.408000000e-07 V_hig
+ 2.408010000e-07 V_hig
+ 2.409000000e-07 V_hig
+ 2.409010000e-07 V_hig
+ 2.410000000e-07 V_hig
+ 2.410010000e-07 V_hig
+ 2.411000000e-07 V_hig
+ 2.411010000e-07 V_hig
+ 2.412000000e-07 V_hig
+ 2.412010000e-07 V_hig
+ 2.413000000e-07 V_hig
+ 2.413010000e-07 V_hig
+ 2.414000000e-07 V_hig
+ 2.414010000e-07 V_hig
+ 2.415000000e-07 V_hig
+ 2.415010000e-07 V_hig
+ 2.416000000e-07 V_hig
+ 2.416010000e-07 V_hig
+ 2.417000000e-07 V_hig
+ 2.417010000e-07 V_hig
+ 2.418000000e-07 V_hig
+ 2.418010000e-07 V_hig
+ 2.419000000e-07 V_hig
+ 2.419010000e-07 V_low
+ 2.420000000e-07 V_low
+ 2.420010000e-07 V_low
+ 2.421000000e-07 V_low
+ 2.421010000e-07 V_low
+ 2.422000000e-07 V_low
+ 2.422010000e-07 V_low
+ 2.423000000e-07 V_low
+ 2.423010000e-07 V_low
+ 2.424000000e-07 V_low
+ 2.424010000e-07 V_low
+ 2.425000000e-07 V_low
+ 2.425010000e-07 V_low
+ 2.426000000e-07 V_low
+ 2.426010000e-07 V_low
+ 2.427000000e-07 V_low
+ 2.427010000e-07 V_low
+ 2.428000000e-07 V_low
+ 2.428010000e-07 V_low
+ 2.429000000e-07 V_low
+ 2.429010000e-07 V_low
+ 2.430000000e-07 V_low
+ 2.430010000e-07 V_low
+ 2.431000000e-07 V_low
+ 2.431010000e-07 V_low
+ 2.432000000e-07 V_low
+ 2.432010000e-07 V_low
+ 2.433000000e-07 V_low
+ 2.433010000e-07 V_low
+ 2.434000000e-07 V_low
+ 2.434010000e-07 V_low
+ 2.435000000e-07 V_low
+ 2.435010000e-07 V_low
+ 2.436000000e-07 V_low
+ 2.436010000e-07 V_low
+ 2.437000000e-07 V_low
+ 2.437010000e-07 V_low
+ 2.438000000e-07 V_low
+ 2.438010000e-07 V_low
+ 2.439000000e-07 V_low
+ 2.439010000e-07 V_low
+ 2.440000000e-07 V_low
+ 2.440010000e-07 V_low
+ 2.441000000e-07 V_low
+ 2.441010000e-07 V_low
+ 2.442000000e-07 V_low
+ 2.442010000e-07 V_low
+ 2.443000000e-07 V_low
+ 2.443010000e-07 V_low
+ 2.444000000e-07 V_low
+ 2.444010000e-07 V_low
+ 2.445000000e-07 V_low
+ 2.445010000e-07 V_low
+ 2.446000000e-07 V_low
+ 2.446010000e-07 V_low
+ 2.447000000e-07 V_low
+ 2.447010000e-07 V_low
+ 2.448000000e-07 V_low
+ 2.448010000e-07 V_low
+ 2.449000000e-07 V_low
+ 2.449010000e-07 V_hig
+ 2.450000000e-07 V_hig
+ 2.450010000e-07 V_hig
+ 2.451000000e-07 V_hig
+ 2.451010000e-07 V_hig
+ 2.452000000e-07 V_hig
+ 2.452010000e-07 V_hig
+ 2.453000000e-07 V_hig
+ 2.453010000e-07 V_hig
+ 2.454000000e-07 V_hig
+ 2.454010000e-07 V_hig
+ 2.455000000e-07 V_hig
+ 2.455010000e-07 V_hig
+ 2.456000000e-07 V_hig
+ 2.456010000e-07 V_hig
+ 2.457000000e-07 V_hig
+ 2.457010000e-07 V_hig
+ 2.458000000e-07 V_hig
+ 2.458010000e-07 V_hig
+ 2.459000000e-07 V_hig
+ 2.459010000e-07 V_hig
+ 2.460000000e-07 V_hig
+ 2.460010000e-07 V_hig
+ 2.461000000e-07 V_hig
+ 2.461010000e-07 V_hig
+ 2.462000000e-07 V_hig
+ 2.462010000e-07 V_hig
+ 2.463000000e-07 V_hig
+ 2.463010000e-07 V_hig
+ 2.464000000e-07 V_hig
+ 2.464010000e-07 V_hig
+ 2.465000000e-07 V_hig
+ 2.465010000e-07 V_hig
+ 2.466000000e-07 V_hig
+ 2.466010000e-07 V_hig
+ 2.467000000e-07 V_hig
+ 2.467010000e-07 V_hig
+ 2.468000000e-07 V_hig
+ 2.468010000e-07 V_hig
+ 2.469000000e-07 V_hig
+ 2.469010000e-07 V_hig
+ 2.470000000e-07 V_hig
+ 2.470010000e-07 V_hig
+ 2.471000000e-07 V_hig
+ 2.471010000e-07 V_hig
+ 2.472000000e-07 V_hig
+ 2.472010000e-07 V_hig
+ 2.473000000e-07 V_hig
+ 2.473010000e-07 V_hig
+ 2.474000000e-07 V_hig
+ 2.474010000e-07 V_hig
+ 2.475000000e-07 V_hig
+ 2.475010000e-07 V_hig
+ 2.476000000e-07 V_hig
+ 2.476010000e-07 V_hig
+ 2.477000000e-07 V_hig
+ 2.477010000e-07 V_hig
+ 2.478000000e-07 V_hig
+ 2.478010000e-07 V_hig
+ 2.479000000e-07 V_hig
+ 2.479010000e-07 V_low
+ 2.480000000e-07 V_low
+ 2.480010000e-07 V_low
+ 2.481000000e-07 V_low
+ 2.481010000e-07 V_low
+ 2.482000000e-07 V_low
+ 2.482010000e-07 V_low
+ 2.483000000e-07 V_low
+ 2.483010000e-07 V_low
+ 2.484000000e-07 V_low
+ 2.484010000e-07 V_low
+ 2.485000000e-07 V_low
+ 2.485010000e-07 V_low
+ 2.486000000e-07 V_low
+ 2.486010000e-07 V_low
+ 2.487000000e-07 V_low
+ 2.487010000e-07 V_low
+ 2.488000000e-07 V_low
+ 2.488010000e-07 V_low
+ 2.489000000e-07 V_low
+ 2.489010000e-07 V_hig
+ 2.490000000e-07 V_hig
+ 2.490010000e-07 V_hig
+ 2.491000000e-07 V_hig
+ 2.491010000e-07 V_hig
+ 2.492000000e-07 V_hig
+ 2.492010000e-07 V_hig
+ 2.493000000e-07 V_hig
+ 2.493010000e-07 V_hig
+ 2.494000000e-07 V_hig
+ 2.494010000e-07 V_hig
+ 2.495000000e-07 V_hig
+ 2.495010000e-07 V_hig
+ 2.496000000e-07 V_hig
+ 2.496010000e-07 V_hig
+ 2.497000000e-07 V_hig
+ 2.497010000e-07 V_hig
+ 2.498000000e-07 V_hig
+ 2.498010000e-07 V_hig
+ 2.499000000e-07 V_hig
+ 2.499010000e-07 V_hig
+ 2.500000000e-07 V_hig
+ 2.500010000e-07 V_hig
+ 2.501000000e-07 V_hig
+ 2.501010000e-07 V_hig
+ 2.502000000e-07 V_hig
+ 2.502010000e-07 V_hig
+ 2.503000000e-07 V_hig
+ 2.503010000e-07 V_hig
+ 2.504000000e-07 V_hig
+ 2.504010000e-07 V_hig
+ 2.505000000e-07 V_hig
+ 2.505010000e-07 V_hig
+ 2.506000000e-07 V_hig
+ 2.506010000e-07 V_hig
+ 2.507000000e-07 V_hig
+ 2.507010000e-07 V_hig
+ 2.508000000e-07 V_hig
+ 2.508010000e-07 V_hig
+ 2.509000000e-07 V_hig
+ 2.509010000e-07 V_low
+ 2.510000000e-07 V_low
+ 2.510010000e-07 V_low
+ 2.511000000e-07 V_low
+ 2.511010000e-07 V_low
+ 2.512000000e-07 V_low
+ 2.512010000e-07 V_low
+ 2.513000000e-07 V_low
+ 2.513010000e-07 V_low
+ 2.514000000e-07 V_low
+ 2.514010000e-07 V_low
+ 2.515000000e-07 V_low
+ 2.515010000e-07 V_low
+ 2.516000000e-07 V_low
+ 2.516010000e-07 V_low
+ 2.517000000e-07 V_low
+ 2.517010000e-07 V_low
+ 2.518000000e-07 V_low
+ 2.518010000e-07 V_low
+ 2.519000000e-07 V_low
+ 2.519010000e-07 V_hig
+ 2.520000000e-07 V_hig
+ 2.520010000e-07 V_hig
+ 2.521000000e-07 V_hig
+ 2.521010000e-07 V_hig
+ 2.522000000e-07 V_hig
+ 2.522010000e-07 V_hig
+ 2.523000000e-07 V_hig
+ 2.523010000e-07 V_hig
+ 2.524000000e-07 V_hig
+ 2.524010000e-07 V_hig
+ 2.525000000e-07 V_hig
+ 2.525010000e-07 V_hig
+ 2.526000000e-07 V_hig
+ 2.526010000e-07 V_hig
+ 2.527000000e-07 V_hig
+ 2.527010000e-07 V_hig
+ 2.528000000e-07 V_hig
+ 2.528010000e-07 V_hig
+ 2.529000000e-07 V_hig
+ 2.529010000e-07 V_low
+ 2.530000000e-07 V_low
+ 2.530010000e-07 V_low
+ 2.531000000e-07 V_low
+ 2.531010000e-07 V_low
+ 2.532000000e-07 V_low
+ 2.532010000e-07 V_low
+ 2.533000000e-07 V_low
+ 2.533010000e-07 V_low
+ 2.534000000e-07 V_low
+ 2.534010000e-07 V_low
+ 2.535000000e-07 V_low
+ 2.535010000e-07 V_low
+ 2.536000000e-07 V_low
+ 2.536010000e-07 V_low
+ 2.537000000e-07 V_low
+ 2.537010000e-07 V_low
+ 2.538000000e-07 V_low
+ 2.538010000e-07 V_low
+ 2.539000000e-07 V_low
+ 2.539010000e-07 V_hig
+ 2.540000000e-07 V_hig
+ 2.540010000e-07 V_hig
+ 2.541000000e-07 V_hig
+ 2.541010000e-07 V_hig
+ 2.542000000e-07 V_hig
+ 2.542010000e-07 V_hig
+ 2.543000000e-07 V_hig
+ 2.543010000e-07 V_hig
+ 2.544000000e-07 V_hig
+ 2.544010000e-07 V_hig
+ 2.545000000e-07 V_hig
+ 2.545010000e-07 V_hig
+ 2.546000000e-07 V_hig
+ 2.546010000e-07 V_hig
+ 2.547000000e-07 V_hig
+ 2.547010000e-07 V_hig
+ 2.548000000e-07 V_hig
+ 2.548010000e-07 V_hig
+ 2.549000000e-07 V_hig
+ 2.549010000e-07 V_hig
+ 2.550000000e-07 V_hig
+ 2.550010000e-07 V_hig
+ 2.551000000e-07 V_hig
+ 2.551010000e-07 V_hig
+ 2.552000000e-07 V_hig
+ 2.552010000e-07 V_hig
+ 2.553000000e-07 V_hig
+ 2.553010000e-07 V_hig
+ 2.554000000e-07 V_hig
+ 2.554010000e-07 V_hig
+ 2.555000000e-07 V_hig
+ 2.555010000e-07 V_hig
+ 2.556000000e-07 V_hig
+ 2.556010000e-07 V_hig
+ 2.557000000e-07 V_hig
+ 2.557010000e-07 V_hig
+ 2.558000000e-07 V_hig
+ 2.558010000e-07 V_hig
+ 2.559000000e-07 V_hig
+ 2.559010000e-07 V_hig
+ 2.560000000e-07 V_hig
+ 2.560010000e-07 V_hig
+ 2.561000000e-07 V_hig
+ 2.561010000e-07 V_hig
+ 2.562000000e-07 V_hig
+ 2.562010000e-07 V_hig
+ 2.563000000e-07 V_hig
+ 2.563010000e-07 V_hig
+ 2.564000000e-07 V_hig
+ 2.564010000e-07 V_hig
+ 2.565000000e-07 V_hig
+ 2.565010000e-07 V_hig
+ 2.566000000e-07 V_hig
+ 2.566010000e-07 V_hig
+ 2.567000000e-07 V_hig
+ 2.567010000e-07 V_hig
+ 2.568000000e-07 V_hig
+ 2.568010000e-07 V_hig
+ 2.569000000e-07 V_hig
+ 2.569010000e-07 V_hig
+ 2.570000000e-07 V_hig
+ 2.570010000e-07 V_hig
+ 2.571000000e-07 V_hig
+ 2.571010000e-07 V_hig
+ 2.572000000e-07 V_hig
+ 2.572010000e-07 V_hig
+ 2.573000000e-07 V_hig
+ 2.573010000e-07 V_hig
+ 2.574000000e-07 V_hig
+ 2.574010000e-07 V_hig
+ 2.575000000e-07 V_hig
+ 2.575010000e-07 V_hig
+ 2.576000000e-07 V_hig
+ 2.576010000e-07 V_hig
+ 2.577000000e-07 V_hig
+ 2.577010000e-07 V_hig
+ 2.578000000e-07 V_hig
+ 2.578010000e-07 V_hig
+ 2.579000000e-07 V_hig
+ 2.579010000e-07 V_low
+ 2.580000000e-07 V_low
+ 2.580010000e-07 V_low
+ 2.581000000e-07 V_low
+ 2.581010000e-07 V_low
+ 2.582000000e-07 V_low
+ 2.582010000e-07 V_low
+ 2.583000000e-07 V_low
+ 2.583010000e-07 V_low
+ 2.584000000e-07 V_low
+ 2.584010000e-07 V_low
+ 2.585000000e-07 V_low
+ 2.585010000e-07 V_low
+ 2.586000000e-07 V_low
+ 2.586010000e-07 V_low
+ 2.587000000e-07 V_low
+ 2.587010000e-07 V_low
+ 2.588000000e-07 V_low
+ 2.588010000e-07 V_low
+ 2.589000000e-07 V_low
+ 2.589010000e-07 V_hig
+ 2.590000000e-07 V_hig
+ 2.590010000e-07 V_hig
+ 2.591000000e-07 V_hig
+ 2.591010000e-07 V_hig
+ 2.592000000e-07 V_hig
+ 2.592010000e-07 V_hig
+ 2.593000000e-07 V_hig
+ 2.593010000e-07 V_hig
+ 2.594000000e-07 V_hig
+ 2.594010000e-07 V_hig
+ 2.595000000e-07 V_hig
+ 2.595010000e-07 V_hig
+ 2.596000000e-07 V_hig
+ 2.596010000e-07 V_hig
+ 2.597000000e-07 V_hig
+ 2.597010000e-07 V_hig
+ 2.598000000e-07 V_hig
+ 2.598010000e-07 V_hig
+ 2.599000000e-07 V_hig
+ 2.599010000e-07 V_low
+ 2.600000000e-07 V_low
+ 2.600010000e-07 V_low
+ 2.601000000e-07 V_low
+ 2.601010000e-07 V_low
+ 2.602000000e-07 V_low
+ 2.602010000e-07 V_low
+ 2.603000000e-07 V_low
+ 2.603010000e-07 V_low
+ 2.604000000e-07 V_low
+ 2.604010000e-07 V_low
+ 2.605000000e-07 V_low
+ 2.605010000e-07 V_low
+ 2.606000000e-07 V_low
+ 2.606010000e-07 V_low
+ 2.607000000e-07 V_low
+ 2.607010000e-07 V_low
+ 2.608000000e-07 V_low
+ 2.608010000e-07 V_low
+ 2.609000000e-07 V_low
+ 2.609010000e-07 V_low
+ 2.610000000e-07 V_low
+ 2.610010000e-07 V_low
+ 2.611000000e-07 V_low
+ 2.611010000e-07 V_low
+ 2.612000000e-07 V_low
+ 2.612010000e-07 V_low
+ 2.613000000e-07 V_low
+ 2.613010000e-07 V_low
+ 2.614000000e-07 V_low
+ 2.614010000e-07 V_low
+ 2.615000000e-07 V_low
+ 2.615010000e-07 V_low
+ 2.616000000e-07 V_low
+ 2.616010000e-07 V_low
+ 2.617000000e-07 V_low
+ 2.617010000e-07 V_low
+ 2.618000000e-07 V_low
+ 2.618010000e-07 V_low
+ 2.619000000e-07 V_low
+ 2.619010000e-07 V_low
+ 2.620000000e-07 V_low
+ 2.620010000e-07 V_low
+ 2.621000000e-07 V_low
+ 2.621010000e-07 V_low
+ 2.622000000e-07 V_low
+ 2.622010000e-07 V_low
+ 2.623000000e-07 V_low
+ 2.623010000e-07 V_low
+ 2.624000000e-07 V_low
+ 2.624010000e-07 V_low
+ 2.625000000e-07 V_low
+ 2.625010000e-07 V_low
+ 2.626000000e-07 V_low
+ 2.626010000e-07 V_low
+ 2.627000000e-07 V_low
+ 2.627010000e-07 V_low
+ 2.628000000e-07 V_low
+ 2.628010000e-07 V_low
+ 2.629000000e-07 V_low
+ 2.629010000e-07 V_hig
+ 2.630000000e-07 V_hig
+ 2.630010000e-07 V_hig
+ 2.631000000e-07 V_hig
+ 2.631010000e-07 V_hig
+ 2.632000000e-07 V_hig
+ 2.632010000e-07 V_hig
+ 2.633000000e-07 V_hig
+ 2.633010000e-07 V_hig
+ 2.634000000e-07 V_hig
+ 2.634010000e-07 V_hig
+ 2.635000000e-07 V_hig
+ 2.635010000e-07 V_hig
+ 2.636000000e-07 V_hig
+ 2.636010000e-07 V_hig
+ 2.637000000e-07 V_hig
+ 2.637010000e-07 V_hig
+ 2.638000000e-07 V_hig
+ 2.638010000e-07 V_hig
+ 2.639000000e-07 V_hig
+ 2.639010000e-07 V_low
+ 2.640000000e-07 V_low
+ 2.640010000e-07 V_low
+ 2.641000000e-07 V_low
+ 2.641010000e-07 V_low
+ 2.642000000e-07 V_low
+ 2.642010000e-07 V_low
+ 2.643000000e-07 V_low
+ 2.643010000e-07 V_low
+ 2.644000000e-07 V_low
+ 2.644010000e-07 V_low
+ 2.645000000e-07 V_low
+ 2.645010000e-07 V_low
+ 2.646000000e-07 V_low
+ 2.646010000e-07 V_low
+ 2.647000000e-07 V_low
+ 2.647010000e-07 V_low
+ 2.648000000e-07 V_low
+ 2.648010000e-07 V_low
+ 2.649000000e-07 V_low
+ 2.649010000e-07 V_low
+ 2.650000000e-07 V_low
+ 2.650010000e-07 V_low
+ 2.651000000e-07 V_low
+ 2.651010000e-07 V_low
+ 2.652000000e-07 V_low
+ 2.652010000e-07 V_low
+ 2.653000000e-07 V_low
+ 2.653010000e-07 V_low
+ 2.654000000e-07 V_low
+ 2.654010000e-07 V_low
+ 2.655000000e-07 V_low
+ 2.655010000e-07 V_low
+ 2.656000000e-07 V_low
+ 2.656010000e-07 V_low
+ 2.657000000e-07 V_low
+ 2.657010000e-07 V_low
+ 2.658000000e-07 V_low
+ 2.658010000e-07 V_low
+ 2.659000000e-07 V_low
+ 2.659010000e-07 V_hig
+ 2.660000000e-07 V_hig
+ 2.660010000e-07 V_hig
+ 2.661000000e-07 V_hig
+ 2.661010000e-07 V_hig
+ 2.662000000e-07 V_hig
+ 2.662010000e-07 V_hig
+ 2.663000000e-07 V_hig
+ 2.663010000e-07 V_hig
+ 2.664000000e-07 V_hig
+ 2.664010000e-07 V_hig
+ 2.665000000e-07 V_hig
+ 2.665010000e-07 V_hig
+ 2.666000000e-07 V_hig
+ 2.666010000e-07 V_hig
+ 2.667000000e-07 V_hig
+ 2.667010000e-07 V_hig
+ 2.668000000e-07 V_hig
+ 2.668010000e-07 V_hig
+ 2.669000000e-07 V_hig
+ 2.669010000e-07 V_hig
+ 2.670000000e-07 V_hig
+ 2.670010000e-07 V_hig
+ 2.671000000e-07 V_hig
+ 2.671010000e-07 V_hig
+ 2.672000000e-07 V_hig
+ 2.672010000e-07 V_hig
+ 2.673000000e-07 V_hig
+ 2.673010000e-07 V_hig
+ 2.674000000e-07 V_hig
+ 2.674010000e-07 V_hig
+ 2.675000000e-07 V_hig
+ 2.675010000e-07 V_hig
+ 2.676000000e-07 V_hig
+ 2.676010000e-07 V_hig
+ 2.677000000e-07 V_hig
+ 2.677010000e-07 V_hig
+ 2.678000000e-07 V_hig
+ 2.678010000e-07 V_hig
+ 2.679000000e-07 V_hig
+ 2.679010000e-07 V_hig
+ 2.680000000e-07 V_hig
+ 2.680010000e-07 V_hig
+ 2.681000000e-07 V_hig
+ 2.681010000e-07 V_hig
+ 2.682000000e-07 V_hig
+ 2.682010000e-07 V_hig
+ 2.683000000e-07 V_hig
+ 2.683010000e-07 V_hig
+ 2.684000000e-07 V_hig
+ 2.684010000e-07 V_hig
+ 2.685000000e-07 V_hig
+ 2.685010000e-07 V_hig
+ 2.686000000e-07 V_hig
+ 2.686010000e-07 V_hig
+ 2.687000000e-07 V_hig
+ 2.687010000e-07 V_hig
+ 2.688000000e-07 V_hig
+ 2.688010000e-07 V_hig
+ 2.689000000e-07 V_hig
+ 2.689010000e-07 V_hig
+ 2.690000000e-07 V_hig
+ 2.690010000e-07 V_hig
+ 2.691000000e-07 V_hig
+ 2.691010000e-07 V_hig
+ 2.692000000e-07 V_hig
+ 2.692010000e-07 V_hig
+ 2.693000000e-07 V_hig
+ 2.693010000e-07 V_hig
+ 2.694000000e-07 V_hig
+ 2.694010000e-07 V_hig
+ 2.695000000e-07 V_hig
+ 2.695010000e-07 V_hig
+ 2.696000000e-07 V_hig
+ 2.696010000e-07 V_hig
+ 2.697000000e-07 V_hig
+ 2.697010000e-07 V_hig
+ 2.698000000e-07 V_hig
+ 2.698010000e-07 V_hig
+ 2.699000000e-07 V_hig
+ 2.699010000e-07 V_low
+ 2.700000000e-07 V_low
+ 2.700010000e-07 V_low
+ 2.701000000e-07 V_low
+ 2.701010000e-07 V_low
+ 2.702000000e-07 V_low
+ 2.702010000e-07 V_low
+ 2.703000000e-07 V_low
+ 2.703010000e-07 V_low
+ 2.704000000e-07 V_low
+ 2.704010000e-07 V_low
+ 2.705000000e-07 V_low
+ 2.705010000e-07 V_low
+ 2.706000000e-07 V_low
+ 2.706010000e-07 V_low
+ 2.707000000e-07 V_low
+ 2.707010000e-07 V_low
+ 2.708000000e-07 V_low
+ 2.708010000e-07 V_low
+ 2.709000000e-07 V_low
+ 2.709010000e-07 V_low
+ 2.710000000e-07 V_low
+ 2.710010000e-07 V_low
+ 2.711000000e-07 V_low
+ 2.711010000e-07 V_low
+ 2.712000000e-07 V_low
+ 2.712010000e-07 V_low
+ 2.713000000e-07 V_low
+ 2.713010000e-07 V_low
+ 2.714000000e-07 V_low
+ 2.714010000e-07 V_low
+ 2.715000000e-07 V_low
+ 2.715010000e-07 V_low
+ 2.716000000e-07 V_low
+ 2.716010000e-07 V_low
+ 2.717000000e-07 V_low
+ 2.717010000e-07 V_low
+ 2.718000000e-07 V_low
+ 2.718010000e-07 V_low
+ 2.719000000e-07 V_low
+ 2.719010000e-07 V_low
+ 2.720000000e-07 V_low
+ 2.720010000e-07 V_low
+ 2.721000000e-07 V_low
+ 2.721010000e-07 V_low
+ 2.722000000e-07 V_low
+ 2.722010000e-07 V_low
+ 2.723000000e-07 V_low
+ 2.723010000e-07 V_low
+ 2.724000000e-07 V_low
+ 2.724010000e-07 V_low
+ 2.725000000e-07 V_low
+ 2.725010000e-07 V_low
+ 2.726000000e-07 V_low
+ 2.726010000e-07 V_low
+ 2.727000000e-07 V_low
+ 2.727010000e-07 V_low
+ 2.728000000e-07 V_low
+ 2.728010000e-07 V_low
+ 2.729000000e-07 V_low
+ 2.729010000e-07 V_hig
+ 2.730000000e-07 V_hig
+ 2.730010000e-07 V_hig
+ 2.731000000e-07 V_hig
+ 2.731010000e-07 V_hig
+ 2.732000000e-07 V_hig
+ 2.732010000e-07 V_hig
+ 2.733000000e-07 V_hig
+ 2.733010000e-07 V_hig
+ 2.734000000e-07 V_hig
+ 2.734010000e-07 V_hig
+ 2.735000000e-07 V_hig
+ 2.735010000e-07 V_hig
+ 2.736000000e-07 V_hig
+ 2.736010000e-07 V_hig
+ 2.737000000e-07 V_hig
+ 2.737010000e-07 V_hig
+ 2.738000000e-07 V_hig
+ 2.738010000e-07 V_hig
+ 2.739000000e-07 V_hig
+ 2.739010000e-07 V_low
+ 2.740000000e-07 V_low
+ 2.740010000e-07 V_low
+ 2.741000000e-07 V_low
+ 2.741010000e-07 V_low
+ 2.742000000e-07 V_low
+ 2.742010000e-07 V_low
+ 2.743000000e-07 V_low
+ 2.743010000e-07 V_low
+ 2.744000000e-07 V_low
+ 2.744010000e-07 V_low
+ 2.745000000e-07 V_low
+ 2.745010000e-07 V_low
+ 2.746000000e-07 V_low
+ 2.746010000e-07 V_low
+ 2.747000000e-07 V_low
+ 2.747010000e-07 V_low
+ 2.748000000e-07 V_low
+ 2.748010000e-07 V_low
+ 2.749000000e-07 V_low
+ 2.749010000e-07 V_low
+ 2.750000000e-07 V_low
+ 2.750010000e-07 V_low
+ 2.751000000e-07 V_low
+ 2.751010000e-07 V_low
+ 2.752000000e-07 V_low
+ 2.752010000e-07 V_low
+ 2.753000000e-07 V_low
+ 2.753010000e-07 V_low
+ 2.754000000e-07 V_low
+ 2.754010000e-07 V_low
+ 2.755000000e-07 V_low
+ 2.755010000e-07 V_low
+ 2.756000000e-07 V_low
+ 2.756010000e-07 V_low
+ 2.757000000e-07 V_low
+ 2.757010000e-07 V_low
+ 2.758000000e-07 V_low
+ 2.758010000e-07 V_low
+ 2.759000000e-07 V_low
+ 2.759010000e-07 V_hig
+ 2.760000000e-07 V_hig
+ 2.760010000e-07 V_hig
+ 2.761000000e-07 V_hig
+ 2.761010000e-07 V_hig
+ 2.762000000e-07 V_hig
+ 2.762010000e-07 V_hig
+ 2.763000000e-07 V_hig
+ 2.763010000e-07 V_hig
+ 2.764000000e-07 V_hig
+ 2.764010000e-07 V_hig
+ 2.765000000e-07 V_hig
+ 2.765010000e-07 V_hig
+ 2.766000000e-07 V_hig
+ 2.766010000e-07 V_hig
+ 2.767000000e-07 V_hig
+ 2.767010000e-07 V_hig
+ 2.768000000e-07 V_hig
+ 2.768010000e-07 V_hig
+ 2.769000000e-07 V_hig
+ 2.769010000e-07 V_hig
+ 2.770000000e-07 V_hig
+ 2.770010000e-07 V_hig
+ 2.771000000e-07 V_hig
+ 2.771010000e-07 V_hig
+ 2.772000000e-07 V_hig
+ 2.772010000e-07 V_hig
+ 2.773000000e-07 V_hig
+ 2.773010000e-07 V_hig
+ 2.774000000e-07 V_hig
+ 2.774010000e-07 V_hig
+ 2.775000000e-07 V_hig
+ 2.775010000e-07 V_hig
+ 2.776000000e-07 V_hig
+ 2.776010000e-07 V_hig
+ 2.777000000e-07 V_hig
+ 2.777010000e-07 V_hig
+ 2.778000000e-07 V_hig
+ 2.778010000e-07 V_hig
+ 2.779000000e-07 V_hig
+ 2.779010000e-07 V_low
+ 2.780000000e-07 V_low
+ 2.780010000e-07 V_low
+ 2.781000000e-07 V_low
+ 2.781010000e-07 V_low
+ 2.782000000e-07 V_low
+ 2.782010000e-07 V_low
+ 2.783000000e-07 V_low
+ 2.783010000e-07 V_low
+ 2.784000000e-07 V_low
+ 2.784010000e-07 V_low
+ 2.785000000e-07 V_low
+ 2.785010000e-07 V_low
+ 2.786000000e-07 V_low
+ 2.786010000e-07 V_low
+ 2.787000000e-07 V_low
+ 2.787010000e-07 V_low
+ 2.788000000e-07 V_low
+ 2.788010000e-07 V_low
+ 2.789000000e-07 V_low
+ 2.789010000e-07 V_low
+ 2.790000000e-07 V_low
+ 2.790010000e-07 V_low
+ 2.791000000e-07 V_low
+ 2.791010000e-07 V_low
+ 2.792000000e-07 V_low
+ 2.792010000e-07 V_low
+ 2.793000000e-07 V_low
+ 2.793010000e-07 V_low
+ 2.794000000e-07 V_low
+ 2.794010000e-07 V_low
+ 2.795000000e-07 V_low
+ 2.795010000e-07 V_low
+ 2.796000000e-07 V_low
+ 2.796010000e-07 V_low
+ 2.797000000e-07 V_low
+ 2.797010000e-07 V_low
+ 2.798000000e-07 V_low
+ 2.798010000e-07 V_low
+ 2.799000000e-07 V_low
+ 2.799010000e-07 V_low
+ 2.800000000e-07 V_low
+ 2.800010000e-07 V_low
+ 2.801000000e-07 V_low
+ 2.801010000e-07 V_low
+ 2.802000000e-07 V_low
+ 2.802010000e-07 V_low
+ 2.803000000e-07 V_low
+ 2.803010000e-07 V_low
+ 2.804000000e-07 V_low
+ 2.804010000e-07 V_low
+ 2.805000000e-07 V_low
+ 2.805010000e-07 V_low
+ 2.806000000e-07 V_low
+ 2.806010000e-07 V_low
+ 2.807000000e-07 V_low
+ 2.807010000e-07 V_low
+ 2.808000000e-07 V_low
+ 2.808010000e-07 V_low
+ 2.809000000e-07 V_low
+ 2.809010000e-07 V_hig
+ 2.810000000e-07 V_hig
+ 2.810010000e-07 V_hig
+ 2.811000000e-07 V_hig
+ 2.811010000e-07 V_hig
+ 2.812000000e-07 V_hig
+ 2.812010000e-07 V_hig
+ 2.813000000e-07 V_hig
+ 2.813010000e-07 V_hig
+ 2.814000000e-07 V_hig
+ 2.814010000e-07 V_hig
+ 2.815000000e-07 V_hig
+ 2.815010000e-07 V_hig
+ 2.816000000e-07 V_hig
+ 2.816010000e-07 V_hig
+ 2.817000000e-07 V_hig
+ 2.817010000e-07 V_hig
+ 2.818000000e-07 V_hig
+ 2.818010000e-07 V_hig
+ 2.819000000e-07 V_hig
+ 2.819010000e-07 V_hig
+ 2.820000000e-07 V_hig
+ 2.820010000e-07 V_hig
+ 2.821000000e-07 V_hig
+ 2.821010000e-07 V_hig
+ 2.822000000e-07 V_hig
+ 2.822010000e-07 V_hig
+ 2.823000000e-07 V_hig
+ 2.823010000e-07 V_hig
+ 2.824000000e-07 V_hig
+ 2.824010000e-07 V_hig
+ 2.825000000e-07 V_hig
+ 2.825010000e-07 V_hig
+ 2.826000000e-07 V_hig
+ 2.826010000e-07 V_hig
+ 2.827000000e-07 V_hig
+ 2.827010000e-07 V_hig
+ 2.828000000e-07 V_hig
+ 2.828010000e-07 V_hig
+ 2.829000000e-07 V_hig
+ 2.829010000e-07 V_hig
+ 2.830000000e-07 V_hig
+ 2.830010000e-07 V_hig
+ 2.831000000e-07 V_hig
+ 2.831010000e-07 V_hig
+ 2.832000000e-07 V_hig
+ 2.832010000e-07 V_hig
+ 2.833000000e-07 V_hig
+ 2.833010000e-07 V_hig
+ 2.834000000e-07 V_hig
+ 2.834010000e-07 V_hig
+ 2.835000000e-07 V_hig
+ 2.835010000e-07 V_hig
+ 2.836000000e-07 V_hig
+ 2.836010000e-07 V_hig
+ 2.837000000e-07 V_hig
+ 2.837010000e-07 V_hig
+ 2.838000000e-07 V_hig
+ 2.838010000e-07 V_hig
+ 2.839000000e-07 V_hig
+ 2.839010000e-07 V_low
+ 2.840000000e-07 V_low
+ 2.840010000e-07 V_low
+ 2.841000000e-07 V_low
+ 2.841010000e-07 V_low
+ 2.842000000e-07 V_low
+ 2.842010000e-07 V_low
+ 2.843000000e-07 V_low
+ 2.843010000e-07 V_low
+ 2.844000000e-07 V_low
+ 2.844010000e-07 V_low
+ 2.845000000e-07 V_low
+ 2.845010000e-07 V_low
+ 2.846000000e-07 V_low
+ 2.846010000e-07 V_low
+ 2.847000000e-07 V_low
+ 2.847010000e-07 V_low
+ 2.848000000e-07 V_low
+ 2.848010000e-07 V_low
+ 2.849000000e-07 V_low
+ 2.849010000e-07 V_hig
+ 2.850000000e-07 V_hig
+ 2.850010000e-07 V_hig
+ 2.851000000e-07 V_hig
+ 2.851010000e-07 V_hig
+ 2.852000000e-07 V_hig
+ 2.852010000e-07 V_hig
+ 2.853000000e-07 V_hig
+ 2.853010000e-07 V_hig
+ 2.854000000e-07 V_hig
+ 2.854010000e-07 V_hig
+ 2.855000000e-07 V_hig
+ 2.855010000e-07 V_hig
+ 2.856000000e-07 V_hig
+ 2.856010000e-07 V_hig
+ 2.857000000e-07 V_hig
+ 2.857010000e-07 V_hig
+ 2.858000000e-07 V_hig
+ 2.858010000e-07 V_hig
+ 2.859000000e-07 V_hig
+ 2.859010000e-07 V_hig
+ 2.860000000e-07 V_hig
+ 2.860010000e-07 V_hig
+ 2.861000000e-07 V_hig
+ 2.861010000e-07 V_hig
+ 2.862000000e-07 V_hig
+ 2.862010000e-07 V_hig
+ 2.863000000e-07 V_hig
+ 2.863010000e-07 V_hig
+ 2.864000000e-07 V_hig
+ 2.864010000e-07 V_hig
+ 2.865000000e-07 V_hig
+ 2.865010000e-07 V_hig
+ 2.866000000e-07 V_hig
+ 2.866010000e-07 V_hig
+ 2.867000000e-07 V_hig
+ 2.867010000e-07 V_hig
+ 2.868000000e-07 V_hig
+ 2.868010000e-07 V_hig
+ 2.869000000e-07 V_hig
+ 2.869010000e-07 V_low
+ 2.870000000e-07 V_low
+ 2.870010000e-07 V_low
+ 2.871000000e-07 V_low
+ 2.871010000e-07 V_low
+ 2.872000000e-07 V_low
+ 2.872010000e-07 V_low
+ 2.873000000e-07 V_low
+ 2.873010000e-07 V_low
+ 2.874000000e-07 V_low
+ 2.874010000e-07 V_low
+ 2.875000000e-07 V_low
+ 2.875010000e-07 V_low
+ 2.876000000e-07 V_low
+ 2.876010000e-07 V_low
+ 2.877000000e-07 V_low
+ 2.877010000e-07 V_low
+ 2.878000000e-07 V_low
+ 2.878010000e-07 V_low
+ 2.879000000e-07 V_low
+ 2.879010000e-07 V_low
+ 2.880000000e-07 V_low
+ 2.880010000e-07 V_low
+ 2.881000000e-07 V_low
+ 2.881010000e-07 V_low
+ 2.882000000e-07 V_low
+ 2.882010000e-07 V_low
+ 2.883000000e-07 V_low
+ 2.883010000e-07 V_low
+ 2.884000000e-07 V_low
+ 2.884010000e-07 V_low
+ 2.885000000e-07 V_low
+ 2.885010000e-07 V_low
+ 2.886000000e-07 V_low
+ 2.886010000e-07 V_low
+ 2.887000000e-07 V_low
+ 2.887010000e-07 V_low
+ 2.888000000e-07 V_low
+ 2.888010000e-07 V_low
+ 2.889000000e-07 V_low
+ 2.889010000e-07 V_low
+ 2.890000000e-07 V_low
+ 2.890010000e-07 V_low
+ 2.891000000e-07 V_low
+ 2.891010000e-07 V_low
+ 2.892000000e-07 V_low
+ 2.892010000e-07 V_low
+ 2.893000000e-07 V_low
+ 2.893010000e-07 V_low
+ 2.894000000e-07 V_low
+ 2.894010000e-07 V_low
+ 2.895000000e-07 V_low
+ 2.895010000e-07 V_low
+ 2.896000000e-07 V_low
+ 2.896010000e-07 V_low
+ 2.897000000e-07 V_low
+ 2.897010000e-07 V_low
+ 2.898000000e-07 V_low
+ 2.898010000e-07 V_low
+ 2.899000000e-07 V_low
+ 2.899010000e-07 V_low
+ 2.900000000e-07 V_low
+ 2.900010000e-07 V_low
+ 2.901000000e-07 V_low
+ 2.901010000e-07 V_low
+ 2.902000000e-07 V_low
+ 2.902010000e-07 V_low
+ 2.903000000e-07 V_low
+ 2.903010000e-07 V_low
+ 2.904000000e-07 V_low
+ 2.904010000e-07 V_low
+ 2.905000000e-07 V_low
+ 2.905010000e-07 V_low
+ 2.906000000e-07 V_low
+ 2.906010000e-07 V_low
+ 2.907000000e-07 V_low
+ 2.907010000e-07 V_low
+ 2.908000000e-07 V_low
+ 2.908010000e-07 V_low
+ 2.909000000e-07 V_low
+ 2.909010000e-07 V_hig
+ 2.910000000e-07 V_hig
+ 2.910010000e-07 V_hig
+ 2.911000000e-07 V_hig
+ 2.911010000e-07 V_hig
+ 2.912000000e-07 V_hig
+ 2.912010000e-07 V_hig
+ 2.913000000e-07 V_hig
+ 2.913010000e-07 V_hig
+ 2.914000000e-07 V_hig
+ 2.914010000e-07 V_hig
+ 2.915000000e-07 V_hig
+ 2.915010000e-07 V_hig
+ 2.916000000e-07 V_hig
+ 2.916010000e-07 V_hig
+ 2.917000000e-07 V_hig
+ 2.917010000e-07 V_hig
+ 2.918000000e-07 V_hig
+ 2.918010000e-07 V_hig
+ 2.919000000e-07 V_hig
+ 2.919010000e-07 V_hig
+ 2.920000000e-07 V_hig
+ 2.920010000e-07 V_hig
+ 2.921000000e-07 V_hig
+ 2.921010000e-07 V_hig
+ 2.922000000e-07 V_hig
+ 2.922010000e-07 V_hig
+ 2.923000000e-07 V_hig
+ 2.923010000e-07 V_hig
+ 2.924000000e-07 V_hig
+ 2.924010000e-07 V_hig
+ 2.925000000e-07 V_hig
+ 2.925010000e-07 V_hig
+ 2.926000000e-07 V_hig
+ 2.926010000e-07 V_hig
+ 2.927000000e-07 V_hig
+ 2.927010000e-07 V_hig
+ 2.928000000e-07 V_hig
+ 2.928010000e-07 V_hig
+ 2.929000000e-07 V_hig
+ 2.929010000e-07 V_hig
+ 2.930000000e-07 V_hig
+ 2.930010000e-07 V_hig
+ 2.931000000e-07 V_hig
+ 2.931010000e-07 V_hig
+ 2.932000000e-07 V_hig
+ 2.932010000e-07 V_hig
+ 2.933000000e-07 V_hig
+ 2.933010000e-07 V_hig
+ 2.934000000e-07 V_hig
+ 2.934010000e-07 V_hig
+ 2.935000000e-07 V_hig
+ 2.935010000e-07 V_hig
+ 2.936000000e-07 V_hig
+ 2.936010000e-07 V_hig
+ 2.937000000e-07 V_hig
+ 2.937010000e-07 V_hig
+ 2.938000000e-07 V_hig
+ 2.938010000e-07 V_hig
+ 2.939000000e-07 V_hig
+ 2.939010000e-07 V_hig
+ 2.940000000e-07 V_hig
+ 2.940010000e-07 V_hig
+ 2.941000000e-07 V_hig
+ 2.941010000e-07 V_hig
+ 2.942000000e-07 V_hig
+ 2.942010000e-07 V_hig
+ 2.943000000e-07 V_hig
+ 2.943010000e-07 V_hig
+ 2.944000000e-07 V_hig
+ 2.944010000e-07 V_hig
+ 2.945000000e-07 V_hig
+ 2.945010000e-07 V_hig
+ 2.946000000e-07 V_hig
+ 2.946010000e-07 V_hig
+ 2.947000000e-07 V_hig
+ 2.947010000e-07 V_hig
+ 2.948000000e-07 V_hig
+ 2.948010000e-07 V_hig
+ 2.949000000e-07 V_hig
+ 2.949010000e-07 V_hig
+ 2.950000000e-07 V_hig
+ 2.950010000e-07 V_hig
+ 2.951000000e-07 V_hig
+ 2.951010000e-07 V_hig
+ 2.952000000e-07 V_hig
+ 2.952010000e-07 V_hig
+ 2.953000000e-07 V_hig
+ 2.953010000e-07 V_hig
+ 2.954000000e-07 V_hig
+ 2.954010000e-07 V_hig
+ 2.955000000e-07 V_hig
+ 2.955010000e-07 V_hig
+ 2.956000000e-07 V_hig
+ 2.956010000e-07 V_hig
+ 2.957000000e-07 V_hig
+ 2.957010000e-07 V_hig
+ 2.958000000e-07 V_hig
+ 2.958010000e-07 V_hig
+ 2.959000000e-07 V_hig
+ 2.959010000e-07 V_hig
+ 2.960000000e-07 V_hig
+ 2.960010000e-07 V_hig
+ 2.961000000e-07 V_hig
+ 2.961010000e-07 V_hig
+ 2.962000000e-07 V_hig
+ 2.962010000e-07 V_hig
+ 2.963000000e-07 V_hig
+ 2.963010000e-07 V_hig
+ 2.964000000e-07 V_hig
+ 2.964010000e-07 V_hig
+ 2.965000000e-07 V_hig
+ 2.965010000e-07 V_hig
+ 2.966000000e-07 V_hig
+ 2.966010000e-07 V_hig
+ 2.967000000e-07 V_hig
+ 2.967010000e-07 V_hig
+ 2.968000000e-07 V_hig
+ 2.968010000e-07 V_hig
+ 2.969000000e-07 V_hig
+ 2.969010000e-07 V_low
+ 2.970000000e-07 V_low
+ 2.970010000e-07 V_low
+ 2.971000000e-07 V_low
+ 2.971010000e-07 V_low
+ 2.972000000e-07 V_low
+ 2.972010000e-07 V_low
+ 2.973000000e-07 V_low
+ 2.973010000e-07 V_low
+ 2.974000000e-07 V_low
+ 2.974010000e-07 V_low
+ 2.975000000e-07 V_low
+ 2.975010000e-07 V_low
+ 2.976000000e-07 V_low
+ 2.976010000e-07 V_low
+ 2.977000000e-07 V_low
+ 2.977010000e-07 V_low
+ 2.978000000e-07 V_low
+ 2.978010000e-07 V_low
+ 2.979000000e-07 V_low
+ 2.979010000e-07 V_hig
+ 2.980000000e-07 V_hig
+ 2.980010000e-07 V_hig
+ 2.981000000e-07 V_hig
+ 2.981010000e-07 V_hig
+ 2.982000000e-07 V_hig
+ 2.982010000e-07 V_hig
+ 2.983000000e-07 V_hig
+ 2.983010000e-07 V_hig
+ 2.984000000e-07 V_hig
+ 2.984010000e-07 V_hig
+ 2.985000000e-07 V_hig
+ 2.985010000e-07 V_hig
+ 2.986000000e-07 V_hig
+ 2.986010000e-07 V_hig
+ 2.987000000e-07 V_hig
+ 2.987010000e-07 V_hig
+ 2.988000000e-07 V_hig
+ 2.988010000e-07 V_hig
+ 2.989000000e-07 V_hig
+ 2.989010000e-07 V_low
+ 2.990000000e-07 V_low
+ 2.990010000e-07 V_low
+ 2.991000000e-07 V_low
+ 2.991010000e-07 V_low
+ 2.992000000e-07 V_low
+ 2.992010000e-07 V_low
+ 2.993000000e-07 V_low
+ 2.993010000e-07 V_low
+ 2.994000000e-07 V_low
+ 2.994010000e-07 V_low
+ 2.995000000e-07 V_low
+ 2.995010000e-07 V_low
+ 2.996000000e-07 V_low
+ 2.996010000e-07 V_low
+ 2.997000000e-07 V_low
+ 2.997010000e-07 V_low
+ 2.998000000e-07 V_low
+ 2.998010000e-07 V_low
+ 2.999000000e-07 V_low
+ 2.999010000e-07 V_low
+ 3.000000000e-07 V_low
+ 3.000010000e-07 V_low
+ 3.001000000e-07 V_low
+ 3.001010000e-07 V_low
+ 3.002000000e-07 V_low
+ 3.002010000e-07 V_low
+ 3.003000000e-07 V_low
+ 3.003010000e-07 V_low
+ 3.004000000e-07 V_low
+ 3.004010000e-07 V_low
+ 3.005000000e-07 V_low
+ 3.005010000e-07 V_low
+ 3.006000000e-07 V_low
+ 3.006010000e-07 V_low
+ 3.007000000e-07 V_low
+ 3.007010000e-07 V_low
+ 3.008000000e-07 V_low
+ 3.008010000e-07 V_low
+ 3.009000000e-07 V_low
+ 3.009010000e-07 V_hig
+ 3.010000000e-07 V_hig
+ 3.010010000e-07 V_hig
+ 3.011000000e-07 V_hig
+ 3.011010000e-07 V_hig
+ 3.012000000e-07 V_hig
+ 3.012010000e-07 V_hig
+ 3.013000000e-07 V_hig
+ 3.013010000e-07 V_hig
+ 3.014000000e-07 V_hig
+ 3.014010000e-07 V_hig
+ 3.015000000e-07 V_hig
+ 3.015010000e-07 V_hig
+ 3.016000000e-07 V_hig
+ 3.016010000e-07 V_hig
+ 3.017000000e-07 V_hig
+ 3.017010000e-07 V_hig
+ 3.018000000e-07 V_hig
+ 3.018010000e-07 V_hig
+ 3.019000000e-07 V_hig
+ 3.019010000e-07 V_hig
+ 3.020000000e-07 V_hig
+ 3.020010000e-07 V_hig
+ 3.021000000e-07 V_hig
+ 3.021010000e-07 V_hig
+ 3.022000000e-07 V_hig
+ 3.022010000e-07 V_hig
+ 3.023000000e-07 V_hig
+ 3.023010000e-07 V_hig
+ 3.024000000e-07 V_hig
+ 3.024010000e-07 V_hig
+ 3.025000000e-07 V_hig
+ 3.025010000e-07 V_hig
+ 3.026000000e-07 V_hig
+ 3.026010000e-07 V_hig
+ 3.027000000e-07 V_hig
+ 3.027010000e-07 V_hig
+ 3.028000000e-07 V_hig
+ 3.028010000e-07 V_hig
+ 3.029000000e-07 V_hig
+ 3.029010000e-07 V_low
+ 3.030000000e-07 V_low
+ 3.030010000e-07 V_low
+ 3.031000000e-07 V_low
+ 3.031010000e-07 V_low
+ 3.032000000e-07 V_low
+ 3.032010000e-07 V_low
+ 3.033000000e-07 V_low
+ 3.033010000e-07 V_low
+ 3.034000000e-07 V_low
+ 3.034010000e-07 V_low
+ 3.035000000e-07 V_low
+ 3.035010000e-07 V_low
+ 3.036000000e-07 V_low
+ 3.036010000e-07 V_low
+ 3.037000000e-07 V_low
+ 3.037010000e-07 V_low
+ 3.038000000e-07 V_low
+ 3.038010000e-07 V_low
+ 3.039000000e-07 V_low
+ 3.039010000e-07 V_low
+ 3.040000000e-07 V_low
+ 3.040010000e-07 V_low
+ 3.041000000e-07 V_low
+ 3.041010000e-07 V_low
+ 3.042000000e-07 V_low
+ 3.042010000e-07 V_low
+ 3.043000000e-07 V_low
+ 3.043010000e-07 V_low
+ 3.044000000e-07 V_low
+ 3.044010000e-07 V_low
+ 3.045000000e-07 V_low
+ 3.045010000e-07 V_low
+ 3.046000000e-07 V_low
+ 3.046010000e-07 V_low
+ 3.047000000e-07 V_low
+ 3.047010000e-07 V_low
+ 3.048000000e-07 V_low
+ 3.048010000e-07 V_low
+ 3.049000000e-07 V_low
+ 3.049010000e-07 V_low
+ 3.050000000e-07 V_low
+ 3.050010000e-07 V_low
+ 3.051000000e-07 V_low
+ 3.051010000e-07 V_low
+ 3.052000000e-07 V_low
+ 3.052010000e-07 V_low
+ 3.053000000e-07 V_low
+ 3.053010000e-07 V_low
+ 3.054000000e-07 V_low
+ 3.054010000e-07 V_low
+ 3.055000000e-07 V_low
+ 3.055010000e-07 V_low
+ 3.056000000e-07 V_low
+ 3.056010000e-07 V_low
+ 3.057000000e-07 V_low
+ 3.057010000e-07 V_low
+ 3.058000000e-07 V_low
+ 3.058010000e-07 V_low
+ 3.059000000e-07 V_low
+ 3.059010000e-07 V_hig
+ 3.060000000e-07 V_hig
+ 3.060010000e-07 V_hig
+ 3.061000000e-07 V_hig
+ 3.061010000e-07 V_hig
+ 3.062000000e-07 V_hig
+ 3.062010000e-07 V_hig
+ 3.063000000e-07 V_hig
+ 3.063010000e-07 V_hig
+ 3.064000000e-07 V_hig
+ 3.064010000e-07 V_hig
+ 3.065000000e-07 V_hig
+ 3.065010000e-07 V_hig
+ 3.066000000e-07 V_hig
+ 3.066010000e-07 V_hig
+ 3.067000000e-07 V_hig
+ 3.067010000e-07 V_hig
+ 3.068000000e-07 V_hig
+ 3.068010000e-07 V_hig
+ 3.069000000e-07 V_hig
+ 3.069010000e-07 V_hig
+ 3.070000000e-07 V_hig
+ 3.070010000e-07 V_hig
+ 3.071000000e-07 V_hig
+ 3.071010000e-07 V_hig
+ 3.072000000e-07 V_hig
+ 3.072010000e-07 V_hig
+ 3.073000000e-07 V_hig
+ 3.073010000e-07 V_hig
+ 3.074000000e-07 V_hig
+ 3.074010000e-07 V_hig
+ 3.075000000e-07 V_hig
+ 3.075010000e-07 V_hig
+ 3.076000000e-07 V_hig
+ 3.076010000e-07 V_hig
+ 3.077000000e-07 V_hig
+ 3.077010000e-07 V_hig
+ 3.078000000e-07 V_hig
+ 3.078010000e-07 V_hig
+ 3.079000000e-07 V_hig
+ 3.079010000e-07 V_low
+ 3.080000000e-07 V_low
+ 3.080010000e-07 V_low
+ 3.081000000e-07 V_low
+ 3.081010000e-07 V_low
+ 3.082000000e-07 V_low
+ 3.082010000e-07 V_low
+ 3.083000000e-07 V_low
+ 3.083010000e-07 V_low
+ 3.084000000e-07 V_low
+ 3.084010000e-07 V_low
+ 3.085000000e-07 V_low
+ 3.085010000e-07 V_low
+ 3.086000000e-07 V_low
+ 3.086010000e-07 V_low
+ 3.087000000e-07 V_low
+ 3.087010000e-07 V_low
+ 3.088000000e-07 V_low
+ 3.088010000e-07 V_low
+ 3.089000000e-07 V_low
+ 3.089010000e-07 V_low
+ 3.090000000e-07 V_low
+ 3.090010000e-07 V_low
+ 3.091000000e-07 V_low
+ 3.091010000e-07 V_low
+ 3.092000000e-07 V_low
+ 3.092010000e-07 V_low
+ 3.093000000e-07 V_low
+ 3.093010000e-07 V_low
+ 3.094000000e-07 V_low
+ 3.094010000e-07 V_low
+ 3.095000000e-07 V_low
+ 3.095010000e-07 V_low
+ 3.096000000e-07 V_low
+ 3.096010000e-07 V_low
+ 3.097000000e-07 V_low
+ 3.097010000e-07 V_low
+ 3.098000000e-07 V_low
+ 3.098010000e-07 V_low
+ 3.099000000e-07 V_low
+ 3.099010000e-07 V_hig
+ 3.100000000e-07 V_hig
+ 3.100010000e-07 V_hig
+ 3.101000000e-07 V_hig
+ 3.101010000e-07 V_hig
+ 3.102000000e-07 V_hig
+ 3.102010000e-07 V_hig
+ 3.103000000e-07 V_hig
+ 3.103010000e-07 V_hig
+ 3.104000000e-07 V_hig
+ 3.104010000e-07 V_hig
+ 3.105000000e-07 V_hig
+ 3.105010000e-07 V_hig
+ 3.106000000e-07 V_hig
+ 3.106010000e-07 V_hig
+ 3.107000000e-07 V_hig
+ 3.107010000e-07 V_hig
+ 3.108000000e-07 V_hig
+ 3.108010000e-07 V_hig
+ 3.109000000e-07 V_hig
+ 3.109010000e-07 V_low
+ 3.110000000e-07 V_low
+ 3.110010000e-07 V_low
+ 3.111000000e-07 V_low
+ 3.111010000e-07 V_low
+ 3.112000000e-07 V_low
+ 3.112010000e-07 V_low
+ 3.113000000e-07 V_low
+ 3.113010000e-07 V_low
+ 3.114000000e-07 V_low
+ 3.114010000e-07 V_low
+ 3.115000000e-07 V_low
+ 3.115010000e-07 V_low
+ 3.116000000e-07 V_low
+ 3.116010000e-07 V_low
+ 3.117000000e-07 V_low
+ 3.117010000e-07 V_low
+ 3.118000000e-07 V_low
+ 3.118010000e-07 V_low
+ 3.119000000e-07 V_low
+ 3.119010000e-07 V_low
+ 3.120000000e-07 V_low
+ 3.120010000e-07 V_low
+ 3.121000000e-07 V_low
+ 3.121010000e-07 V_low
+ 3.122000000e-07 V_low
+ 3.122010000e-07 V_low
+ 3.123000000e-07 V_low
+ 3.123010000e-07 V_low
+ 3.124000000e-07 V_low
+ 3.124010000e-07 V_low
+ 3.125000000e-07 V_low
+ 3.125010000e-07 V_low
+ 3.126000000e-07 V_low
+ 3.126010000e-07 V_low
+ 3.127000000e-07 V_low
+ 3.127010000e-07 V_low
+ 3.128000000e-07 V_low
+ 3.128010000e-07 V_low
+ 3.129000000e-07 V_low
+ 3.129010000e-07 V_low
+ 3.130000000e-07 V_low
+ 3.130010000e-07 V_low
+ 3.131000000e-07 V_low
+ 3.131010000e-07 V_low
+ 3.132000000e-07 V_low
+ 3.132010000e-07 V_low
+ 3.133000000e-07 V_low
+ 3.133010000e-07 V_low
+ 3.134000000e-07 V_low
+ 3.134010000e-07 V_low
+ 3.135000000e-07 V_low
+ 3.135010000e-07 V_low
+ 3.136000000e-07 V_low
+ 3.136010000e-07 V_low
+ 3.137000000e-07 V_low
+ 3.137010000e-07 V_low
+ 3.138000000e-07 V_low
+ 3.138010000e-07 V_low
+ 3.139000000e-07 V_low
+ 3.139010000e-07 V_hig
+ 3.140000000e-07 V_hig
+ 3.140010000e-07 V_hig
+ 3.141000000e-07 V_hig
+ 3.141010000e-07 V_hig
+ 3.142000000e-07 V_hig
+ 3.142010000e-07 V_hig
+ 3.143000000e-07 V_hig
+ 3.143010000e-07 V_hig
+ 3.144000000e-07 V_hig
+ 3.144010000e-07 V_hig
+ 3.145000000e-07 V_hig
+ 3.145010000e-07 V_hig
+ 3.146000000e-07 V_hig
+ 3.146010000e-07 V_hig
+ 3.147000000e-07 V_hig
+ 3.147010000e-07 V_hig
+ 3.148000000e-07 V_hig
+ 3.148010000e-07 V_hig
+ 3.149000000e-07 V_hig
+ 3.149010000e-07 V_low
+ 3.150000000e-07 V_low
+ 3.150010000e-07 V_low
+ 3.151000000e-07 V_low
+ 3.151010000e-07 V_low
+ 3.152000000e-07 V_low
+ 3.152010000e-07 V_low
+ 3.153000000e-07 V_low
+ 3.153010000e-07 V_low
+ 3.154000000e-07 V_low
+ 3.154010000e-07 V_low
+ 3.155000000e-07 V_low
+ 3.155010000e-07 V_low
+ 3.156000000e-07 V_low
+ 3.156010000e-07 V_low
+ 3.157000000e-07 V_low
+ 3.157010000e-07 V_low
+ 3.158000000e-07 V_low
+ 3.158010000e-07 V_low
+ 3.159000000e-07 V_low
+ 3.159010000e-07 V_low
+ 3.160000000e-07 V_low
+ 3.160010000e-07 V_low
+ 3.161000000e-07 V_low
+ 3.161010000e-07 V_low
+ 3.162000000e-07 V_low
+ 3.162010000e-07 V_low
+ 3.163000000e-07 V_low
+ 3.163010000e-07 V_low
+ 3.164000000e-07 V_low
+ 3.164010000e-07 V_low
+ 3.165000000e-07 V_low
+ 3.165010000e-07 V_low
+ 3.166000000e-07 V_low
+ 3.166010000e-07 V_low
+ 3.167000000e-07 V_low
+ 3.167010000e-07 V_low
+ 3.168000000e-07 V_low
+ 3.168010000e-07 V_low
+ 3.169000000e-07 V_low
+ 3.169010000e-07 V_low
+ 3.170000000e-07 V_low
+ 3.170010000e-07 V_low
+ 3.171000000e-07 V_low
+ 3.171010000e-07 V_low
+ 3.172000000e-07 V_low
+ 3.172010000e-07 V_low
+ 3.173000000e-07 V_low
+ 3.173010000e-07 V_low
+ 3.174000000e-07 V_low
+ 3.174010000e-07 V_low
+ 3.175000000e-07 V_low
+ 3.175010000e-07 V_low
+ 3.176000000e-07 V_low
+ 3.176010000e-07 V_low
+ 3.177000000e-07 V_low
+ 3.177010000e-07 V_low
+ 3.178000000e-07 V_low
+ 3.178010000e-07 V_low
+ 3.179000000e-07 V_low
+ 3.179010000e-07 V_hig
+ 3.180000000e-07 V_hig
+ 3.180010000e-07 V_hig
+ 3.181000000e-07 V_hig
+ 3.181010000e-07 V_hig
+ 3.182000000e-07 V_hig
+ 3.182010000e-07 V_hig
+ 3.183000000e-07 V_hig
+ 3.183010000e-07 V_hig
+ 3.184000000e-07 V_hig
+ 3.184010000e-07 V_hig
+ 3.185000000e-07 V_hig
+ 3.185010000e-07 V_hig
+ 3.186000000e-07 V_hig
+ 3.186010000e-07 V_hig
+ 3.187000000e-07 V_hig
+ 3.187010000e-07 V_hig
+ 3.188000000e-07 V_hig
+ 3.188010000e-07 V_hig
+ 3.189000000e-07 V_hig
+ 3.189010000e-07 V_low
+ 3.190000000e-07 V_low
+ 3.190010000e-07 V_low
+ 3.191000000e-07 V_low
+ 3.191010000e-07 V_low
+ 3.192000000e-07 V_low
+ 3.192010000e-07 V_low
+ 3.193000000e-07 V_low
+ 3.193010000e-07 V_low
+ 3.194000000e-07 V_low
+ 3.194010000e-07 V_low
+ 3.195000000e-07 V_low
+ 3.195010000e-07 V_low
+ 3.196000000e-07 V_low
+ 3.196010000e-07 V_low
+ 3.197000000e-07 V_low
+ 3.197010000e-07 V_low
+ 3.198000000e-07 V_low
+ 3.198010000e-07 V_low
+ 3.199000000e-07 V_low
+ 3.199010000e-07 V_hig
+ 3.200000000e-07 V_hig
+ 3.200010000e-07 V_hig
+ 3.201000000e-07 V_hig
+ 3.201010000e-07 V_hig
+ 3.202000000e-07 V_hig
+ 3.202010000e-07 V_hig
+ 3.203000000e-07 V_hig
+ 3.203010000e-07 V_hig
+ 3.204000000e-07 V_hig
+ 3.204010000e-07 V_hig
+ 3.205000000e-07 V_hig
+ 3.205010000e-07 V_hig
+ 3.206000000e-07 V_hig
+ 3.206010000e-07 V_hig
+ 3.207000000e-07 V_hig
+ 3.207010000e-07 V_hig
+ 3.208000000e-07 V_hig
+ 3.208010000e-07 V_hig
+ 3.209000000e-07 V_hig
+ 3.209010000e-07 V_low
+ 3.210000000e-07 V_low
+ 3.210010000e-07 V_low
+ 3.211000000e-07 V_low
+ 3.211010000e-07 V_low
+ 3.212000000e-07 V_low
+ 3.212010000e-07 V_low
+ 3.213000000e-07 V_low
+ 3.213010000e-07 V_low
+ 3.214000000e-07 V_low
+ 3.214010000e-07 V_low
+ 3.215000000e-07 V_low
+ 3.215010000e-07 V_low
+ 3.216000000e-07 V_low
+ 3.216010000e-07 V_low
+ 3.217000000e-07 V_low
+ 3.217010000e-07 V_low
+ 3.218000000e-07 V_low
+ 3.218010000e-07 V_low
+ 3.219000000e-07 V_low
+ 3.219010000e-07 V_hig
+ 3.220000000e-07 V_hig
+ 3.220010000e-07 V_hig
+ 3.221000000e-07 V_hig
+ 3.221010000e-07 V_hig
+ 3.222000000e-07 V_hig
+ 3.222010000e-07 V_hig
+ 3.223000000e-07 V_hig
+ 3.223010000e-07 V_hig
+ 3.224000000e-07 V_hig
+ 3.224010000e-07 V_hig
+ 3.225000000e-07 V_hig
+ 3.225010000e-07 V_hig
+ 3.226000000e-07 V_hig
+ 3.226010000e-07 V_hig
+ 3.227000000e-07 V_hig
+ 3.227010000e-07 V_hig
+ 3.228000000e-07 V_hig
+ 3.228010000e-07 V_hig
+ 3.229000000e-07 V_hig
+ 3.229010000e-07 V_low
+ 3.230000000e-07 V_low
+ 3.230010000e-07 V_low
+ 3.231000000e-07 V_low
+ 3.231010000e-07 V_low
+ 3.232000000e-07 V_low
+ 3.232010000e-07 V_low
+ 3.233000000e-07 V_low
+ 3.233010000e-07 V_low
+ 3.234000000e-07 V_low
+ 3.234010000e-07 V_low
+ 3.235000000e-07 V_low
+ 3.235010000e-07 V_low
+ 3.236000000e-07 V_low
+ 3.236010000e-07 V_low
+ 3.237000000e-07 V_low
+ 3.237010000e-07 V_low
+ 3.238000000e-07 V_low
+ 3.238010000e-07 V_low
+ 3.239000000e-07 V_low
+ 3.239010000e-07 V_low
+ 3.240000000e-07 V_low
+ 3.240010000e-07 V_low
+ 3.241000000e-07 V_low
+ 3.241010000e-07 V_low
+ 3.242000000e-07 V_low
+ 3.242010000e-07 V_low
+ 3.243000000e-07 V_low
+ 3.243010000e-07 V_low
+ 3.244000000e-07 V_low
+ 3.244010000e-07 V_low
+ 3.245000000e-07 V_low
+ 3.245010000e-07 V_low
+ 3.246000000e-07 V_low
+ 3.246010000e-07 V_low
+ 3.247000000e-07 V_low
+ 3.247010000e-07 V_low
+ 3.248000000e-07 V_low
+ 3.248010000e-07 V_low
+ 3.249000000e-07 V_low
+ 3.249010000e-07 V_hig
+ 3.250000000e-07 V_hig
+ 3.250010000e-07 V_hig
+ 3.251000000e-07 V_hig
+ 3.251010000e-07 V_hig
+ 3.252000000e-07 V_hig
+ 3.252010000e-07 V_hig
+ 3.253000000e-07 V_hig
+ 3.253010000e-07 V_hig
+ 3.254000000e-07 V_hig
+ 3.254010000e-07 V_hig
+ 3.255000000e-07 V_hig
+ 3.255010000e-07 V_hig
+ 3.256000000e-07 V_hig
+ 3.256010000e-07 V_hig
+ 3.257000000e-07 V_hig
+ 3.257010000e-07 V_hig
+ 3.258000000e-07 V_hig
+ 3.258010000e-07 V_hig
+ 3.259000000e-07 V_hig
+ 3.259010000e-07 V_low
+ 3.260000000e-07 V_low
+ 3.260010000e-07 V_low
+ 3.261000000e-07 V_low
+ 3.261010000e-07 V_low
+ 3.262000000e-07 V_low
+ 3.262010000e-07 V_low
+ 3.263000000e-07 V_low
+ 3.263010000e-07 V_low
+ 3.264000000e-07 V_low
+ 3.264010000e-07 V_low
+ 3.265000000e-07 V_low
+ 3.265010000e-07 V_low
+ 3.266000000e-07 V_low
+ 3.266010000e-07 V_low
+ 3.267000000e-07 V_low
+ 3.267010000e-07 V_low
+ 3.268000000e-07 V_low
+ 3.268010000e-07 V_low
+ 3.269000000e-07 V_low
+ 3.269010000e-07 V_low
+ 3.270000000e-07 V_low
+ 3.270010000e-07 V_low
+ 3.271000000e-07 V_low
+ 3.271010000e-07 V_low
+ 3.272000000e-07 V_low
+ 3.272010000e-07 V_low
+ 3.273000000e-07 V_low
+ 3.273010000e-07 V_low
+ 3.274000000e-07 V_low
+ 3.274010000e-07 V_low
+ 3.275000000e-07 V_low
+ 3.275010000e-07 V_low
+ 3.276000000e-07 V_low
+ 3.276010000e-07 V_low
+ 3.277000000e-07 V_low
+ 3.277010000e-07 V_low
+ 3.278000000e-07 V_low
+ 3.278010000e-07 V_low
+ 3.279000000e-07 V_low
+ 3.279010000e-07 V_hig
+ 3.280000000e-07 V_hig
+ 3.280010000e-07 V_hig
+ 3.281000000e-07 V_hig
+ 3.281010000e-07 V_hig
+ 3.282000000e-07 V_hig
+ 3.282010000e-07 V_hig
+ 3.283000000e-07 V_hig
+ 3.283010000e-07 V_hig
+ 3.284000000e-07 V_hig
+ 3.284010000e-07 V_hig
+ 3.285000000e-07 V_hig
+ 3.285010000e-07 V_hig
+ 3.286000000e-07 V_hig
+ 3.286010000e-07 V_hig
+ 3.287000000e-07 V_hig
+ 3.287010000e-07 V_hig
+ 3.288000000e-07 V_hig
+ 3.288010000e-07 V_hig
+ 3.289000000e-07 V_hig
+ 3.289010000e-07 V_hig
+ 3.290000000e-07 V_hig
+ 3.290010000e-07 V_hig
+ 3.291000000e-07 V_hig
+ 3.291010000e-07 V_hig
+ 3.292000000e-07 V_hig
+ 3.292010000e-07 V_hig
+ 3.293000000e-07 V_hig
+ 3.293010000e-07 V_hig
+ 3.294000000e-07 V_hig
+ 3.294010000e-07 V_hig
+ 3.295000000e-07 V_hig
+ 3.295010000e-07 V_hig
+ 3.296000000e-07 V_hig
+ 3.296010000e-07 V_hig
+ 3.297000000e-07 V_hig
+ 3.297010000e-07 V_hig
+ 3.298000000e-07 V_hig
+ 3.298010000e-07 V_hig
+ 3.299000000e-07 V_hig
+ 3.299010000e-07 V_hig
+ 3.300000000e-07 V_hig
+ 3.300010000e-07 V_hig
+ 3.301000000e-07 V_hig
+ 3.301010000e-07 V_hig
+ 3.302000000e-07 V_hig
+ 3.302010000e-07 V_hig
+ 3.303000000e-07 V_hig
+ 3.303010000e-07 V_hig
+ 3.304000000e-07 V_hig
+ 3.304010000e-07 V_hig
+ 3.305000000e-07 V_hig
+ 3.305010000e-07 V_hig
+ 3.306000000e-07 V_hig
+ 3.306010000e-07 V_hig
+ 3.307000000e-07 V_hig
+ 3.307010000e-07 V_hig
+ 3.308000000e-07 V_hig
+ 3.308010000e-07 V_hig
+ 3.309000000e-07 V_hig
+ 3.309010000e-07 V_low
+ 3.310000000e-07 V_low
+ 3.310010000e-07 V_low
+ 3.311000000e-07 V_low
+ 3.311010000e-07 V_low
+ 3.312000000e-07 V_low
+ 3.312010000e-07 V_low
+ 3.313000000e-07 V_low
+ 3.313010000e-07 V_low
+ 3.314000000e-07 V_low
+ 3.314010000e-07 V_low
+ 3.315000000e-07 V_low
+ 3.315010000e-07 V_low
+ 3.316000000e-07 V_low
+ 3.316010000e-07 V_low
+ 3.317000000e-07 V_low
+ 3.317010000e-07 V_low
+ 3.318000000e-07 V_low
+ 3.318010000e-07 V_low
+ 3.319000000e-07 V_low
+ 3.319010000e-07 V_hig
+ 3.320000000e-07 V_hig
+ 3.320010000e-07 V_hig
+ 3.321000000e-07 V_hig
+ 3.321010000e-07 V_hig
+ 3.322000000e-07 V_hig
+ 3.322010000e-07 V_hig
+ 3.323000000e-07 V_hig
+ 3.323010000e-07 V_hig
+ 3.324000000e-07 V_hig
+ 3.324010000e-07 V_hig
+ 3.325000000e-07 V_hig
+ 3.325010000e-07 V_hig
+ 3.326000000e-07 V_hig
+ 3.326010000e-07 V_hig
+ 3.327000000e-07 V_hig
+ 3.327010000e-07 V_hig
+ 3.328000000e-07 V_hig
+ 3.328010000e-07 V_hig
+ 3.329000000e-07 V_hig
+ 3.329010000e-07 V_hig
+ 3.330000000e-07 V_hig
+ 3.330010000e-07 V_hig
+ 3.331000000e-07 V_hig
+ 3.331010000e-07 V_hig
+ 3.332000000e-07 V_hig
+ 3.332010000e-07 V_hig
+ 3.333000000e-07 V_hig
+ 3.333010000e-07 V_hig
+ 3.334000000e-07 V_hig
+ 3.334010000e-07 V_hig
+ 3.335000000e-07 V_hig
+ 3.335010000e-07 V_hig
+ 3.336000000e-07 V_hig
+ 3.336010000e-07 V_hig
+ 3.337000000e-07 V_hig
+ 3.337010000e-07 V_hig
+ 3.338000000e-07 V_hig
+ 3.338010000e-07 V_hig
+ 3.339000000e-07 V_hig
+ 3.339010000e-07 V_low
+ 3.340000000e-07 V_low
+ 3.340010000e-07 V_low
+ 3.341000000e-07 V_low
+ 3.341010000e-07 V_low
+ 3.342000000e-07 V_low
+ 3.342010000e-07 V_low
+ 3.343000000e-07 V_low
+ 3.343010000e-07 V_low
+ 3.344000000e-07 V_low
+ 3.344010000e-07 V_low
+ 3.345000000e-07 V_low
+ 3.345010000e-07 V_low
+ 3.346000000e-07 V_low
+ 3.346010000e-07 V_low
+ 3.347000000e-07 V_low
+ 3.347010000e-07 V_low
+ 3.348000000e-07 V_low
+ 3.348010000e-07 V_low
+ 3.349000000e-07 V_low
+ 3.349010000e-07 V_hig
+ 3.350000000e-07 V_hig
+ 3.350010000e-07 V_hig
+ 3.351000000e-07 V_hig
+ 3.351010000e-07 V_hig
+ 3.352000000e-07 V_hig
+ 3.352010000e-07 V_hig
+ 3.353000000e-07 V_hig
+ 3.353010000e-07 V_hig
+ 3.354000000e-07 V_hig
+ 3.354010000e-07 V_hig
+ 3.355000000e-07 V_hig
+ 3.355010000e-07 V_hig
+ 3.356000000e-07 V_hig
+ 3.356010000e-07 V_hig
+ 3.357000000e-07 V_hig
+ 3.357010000e-07 V_hig
+ 3.358000000e-07 V_hig
+ 3.358010000e-07 V_hig
+ 3.359000000e-07 V_hig
+ 3.359010000e-07 V_hig
+ 3.360000000e-07 V_hig
+ 3.360010000e-07 V_hig
+ 3.361000000e-07 V_hig
+ 3.361010000e-07 V_hig
+ 3.362000000e-07 V_hig
+ 3.362010000e-07 V_hig
+ 3.363000000e-07 V_hig
+ 3.363010000e-07 V_hig
+ 3.364000000e-07 V_hig
+ 3.364010000e-07 V_hig
+ 3.365000000e-07 V_hig
+ 3.365010000e-07 V_hig
+ 3.366000000e-07 V_hig
+ 3.366010000e-07 V_hig
+ 3.367000000e-07 V_hig
+ 3.367010000e-07 V_hig
+ 3.368000000e-07 V_hig
+ 3.368010000e-07 V_hig
+ 3.369000000e-07 V_hig
+ 3.369010000e-07 V_low
+ 3.370000000e-07 V_low
+ 3.370010000e-07 V_low
+ 3.371000000e-07 V_low
+ 3.371010000e-07 V_low
+ 3.372000000e-07 V_low
+ 3.372010000e-07 V_low
+ 3.373000000e-07 V_low
+ 3.373010000e-07 V_low
+ 3.374000000e-07 V_low
+ 3.374010000e-07 V_low
+ 3.375000000e-07 V_low
+ 3.375010000e-07 V_low
+ 3.376000000e-07 V_low
+ 3.376010000e-07 V_low
+ 3.377000000e-07 V_low
+ 3.377010000e-07 V_low
+ 3.378000000e-07 V_low
+ 3.378010000e-07 V_low
+ 3.379000000e-07 V_low
+ 3.379010000e-07 V_low
+ 3.380000000e-07 V_low
+ 3.380010000e-07 V_low
+ 3.381000000e-07 V_low
+ 3.381010000e-07 V_low
+ 3.382000000e-07 V_low
+ 3.382010000e-07 V_low
+ 3.383000000e-07 V_low
+ 3.383010000e-07 V_low
+ 3.384000000e-07 V_low
+ 3.384010000e-07 V_low
+ 3.385000000e-07 V_low
+ 3.385010000e-07 V_low
+ 3.386000000e-07 V_low
+ 3.386010000e-07 V_low
+ 3.387000000e-07 V_low
+ 3.387010000e-07 V_low
+ 3.388000000e-07 V_low
+ 3.388010000e-07 V_low
+ 3.389000000e-07 V_low
+ 3.389010000e-07 V_hig
+ 3.390000000e-07 V_hig
+ 3.390010000e-07 V_hig
+ 3.391000000e-07 V_hig
+ 3.391010000e-07 V_hig
+ 3.392000000e-07 V_hig
+ 3.392010000e-07 V_hig
+ 3.393000000e-07 V_hig
+ 3.393010000e-07 V_hig
+ 3.394000000e-07 V_hig
+ 3.394010000e-07 V_hig
+ 3.395000000e-07 V_hig
+ 3.395010000e-07 V_hig
+ 3.396000000e-07 V_hig
+ 3.396010000e-07 V_hig
+ 3.397000000e-07 V_hig
+ 3.397010000e-07 V_hig
+ 3.398000000e-07 V_hig
+ 3.398010000e-07 V_hig
+ 3.399000000e-07 V_hig
+ 3.399010000e-07 V_low
+ 3.400000000e-07 V_low
+ 3.400010000e-07 V_low
+ 3.401000000e-07 V_low
+ 3.401010000e-07 V_low
+ 3.402000000e-07 V_low
+ 3.402010000e-07 V_low
+ 3.403000000e-07 V_low
+ 3.403010000e-07 V_low
+ 3.404000000e-07 V_low
+ 3.404010000e-07 V_low
+ 3.405000000e-07 V_low
+ 3.405010000e-07 V_low
+ 3.406000000e-07 V_low
+ 3.406010000e-07 V_low
+ 3.407000000e-07 V_low
+ 3.407010000e-07 V_low
+ 3.408000000e-07 V_low
+ 3.408010000e-07 V_low
+ 3.409000000e-07 V_low
+ 3.409010000e-07 V_low
+ 3.410000000e-07 V_low
+ 3.410010000e-07 V_low
+ 3.411000000e-07 V_low
+ 3.411010000e-07 V_low
+ 3.412000000e-07 V_low
+ 3.412010000e-07 V_low
+ 3.413000000e-07 V_low
+ 3.413010000e-07 V_low
+ 3.414000000e-07 V_low
+ 3.414010000e-07 V_low
+ 3.415000000e-07 V_low
+ 3.415010000e-07 V_low
+ 3.416000000e-07 V_low
+ 3.416010000e-07 V_low
+ 3.417000000e-07 V_low
+ 3.417010000e-07 V_low
+ 3.418000000e-07 V_low
+ 3.418010000e-07 V_low
+ 3.419000000e-07 V_low
+ 3.419010000e-07 V_low
+ 3.420000000e-07 V_low
+ 3.420010000e-07 V_low
+ 3.421000000e-07 V_low
+ 3.421010000e-07 V_low
+ 3.422000000e-07 V_low
+ 3.422010000e-07 V_low
+ 3.423000000e-07 V_low
+ 3.423010000e-07 V_low
+ 3.424000000e-07 V_low
+ 3.424010000e-07 V_low
+ 3.425000000e-07 V_low
+ 3.425010000e-07 V_low
+ 3.426000000e-07 V_low
+ 3.426010000e-07 V_low
+ 3.427000000e-07 V_low
+ 3.427010000e-07 V_low
+ 3.428000000e-07 V_low
+ 3.428010000e-07 V_low
+ 3.429000000e-07 V_low
+ 3.429010000e-07 V_hig
+ 3.430000000e-07 V_hig
+ 3.430010000e-07 V_hig
+ 3.431000000e-07 V_hig
+ 3.431010000e-07 V_hig
+ 3.432000000e-07 V_hig
+ 3.432010000e-07 V_hig
+ 3.433000000e-07 V_hig
+ 3.433010000e-07 V_hig
+ 3.434000000e-07 V_hig
+ 3.434010000e-07 V_hig
+ 3.435000000e-07 V_hig
+ 3.435010000e-07 V_hig
+ 3.436000000e-07 V_hig
+ 3.436010000e-07 V_hig
+ 3.437000000e-07 V_hig
+ 3.437010000e-07 V_hig
+ 3.438000000e-07 V_hig
+ 3.438010000e-07 V_hig
+ 3.439000000e-07 V_hig
+ 3.439010000e-07 V_hig
+ 3.440000000e-07 V_hig
+ 3.440010000e-07 V_hig
+ 3.441000000e-07 V_hig
+ 3.441010000e-07 V_hig
+ 3.442000000e-07 V_hig
+ 3.442010000e-07 V_hig
+ 3.443000000e-07 V_hig
+ 3.443010000e-07 V_hig
+ 3.444000000e-07 V_hig
+ 3.444010000e-07 V_hig
+ 3.445000000e-07 V_hig
+ 3.445010000e-07 V_hig
+ 3.446000000e-07 V_hig
+ 3.446010000e-07 V_hig
+ 3.447000000e-07 V_hig
+ 3.447010000e-07 V_hig
+ 3.448000000e-07 V_hig
+ 3.448010000e-07 V_hig
+ 3.449000000e-07 V_hig
+ 3.449010000e-07 V_low
+ 3.450000000e-07 V_low
+ 3.450010000e-07 V_low
+ 3.451000000e-07 V_low
+ 3.451010000e-07 V_low
+ 3.452000000e-07 V_low
+ 3.452010000e-07 V_low
+ 3.453000000e-07 V_low
+ 3.453010000e-07 V_low
+ 3.454000000e-07 V_low
+ 3.454010000e-07 V_low
+ 3.455000000e-07 V_low
+ 3.455010000e-07 V_low
+ 3.456000000e-07 V_low
+ 3.456010000e-07 V_low
+ 3.457000000e-07 V_low
+ 3.457010000e-07 V_low
+ 3.458000000e-07 V_low
+ 3.458010000e-07 V_low
+ 3.459000000e-07 V_low
+ 3.459010000e-07 V_low
+ 3.460000000e-07 V_low
+ 3.460010000e-07 V_low
+ 3.461000000e-07 V_low
+ 3.461010000e-07 V_low
+ 3.462000000e-07 V_low
+ 3.462010000e-07 V_low
+ 3.463000000e-07 V_low
+ 3.463010000e-07 V_low
+ 3.464000000e-07 V_low
+ 3.464010000e-07 V_low
+ 3.465000000e-07 V_low
+ 3.465010000e-07 V_low
+ 3.466000000e-07 V_low
+ 3.466010000e-07 V_low
+ 3.467000000e-07 V_low
+ 3.467010000e-07 V_low
+ 3.468000000e-07 V_low
+ 3.468010000e-07 V_low
+ 3.469000000e-07 V_low
+ 3.469010000e-07 V_hig
+ 3.470000000e-07 V_hig
+ 3.470010000e-07 V_hig
+ 3.471000000e-07 V_hig
+ 3.471010000e-07 V_hig
+ 3.472000000e-07 V_hig
+ 3.472010000e-07 V_hig
+ 3.473000000e-07 V_hig
+ 3.473010000e-07 V_hig
+ 3.474000000e-07 V_hig
+ 3.474010000e-07 V_hig
+ 3.475000000e-07 V_hig
+ 3.475010000e-07 V_hig
+ 3.476000000e-07 V_hig
+ 3.476010000e-07 V_hig
+ 3.477000000e-07 V_hig
+ 3.477010000e-07 V_hig
+ 3.478000000e-07 V_hig
+ 3.478010000e-07 V_hig
+ 3.479000000e-07 V_hig
+ 3.479010000e-07 V_low
+ 3.480000000e-07 V_low
+ 3.480010000e-07 V_low
+ 3.481000000e-07 V_low
+ 3.481010000e-07 V_low
+ 3.482000000e-07 V_low
+ 3.482010000e-07 V_low
+ 3.483000000e-07 V_low
+ 3.483010000e-07 V_low
+ 3.484000000e-07 V_low
+ 3.484010000e-07 V_low
+ 3.485000000e-07 V_low
+ 3.485010000e-07 V_low
+ 3.486000000e-07 V_low
+ 3.486010000e-07 V_low
+ 3.487000000e-07 V_low
+ 3.487010000e-07 V_low
+ 3.488000000e-07 V_low
+ 3.488010000e-07 V_low
+ 3.489000000e-07 V_low
+ 3.489010000e-07 V_low
+ 3.490000000e-07 V_low
+ 3.490010000e-07 V_low
+ 3.491000000e-07 V_low
+ 3.491010000e-07 V_low
+ 3.492000000e-07 V_low
+ 3.492010000e-07 V_low
+ 3.493000000e-07 V_low
+ 3.493010000e-07 V_low
+ 3.494000000e-07 V_low
+ 3.494010000e-07 V_low
+ 3.495000000e-07 V_low
+ 3.495010000e-07 V_low
+ 3.496000000e-07 V_low
+ 3.496010000e-07 V_low
+ 3.497000000e-07 V_low
+ 3.497010000e-07 V_low
+ 3.498000000e-07 V_low
+ 3.498010000e-07 V_low
+ 3.499000000e-07 V_low
+ 3.499010000e-07 V_hig
+ 3.500000000e-07 V_hig
+ 3.500010000e-07 V_hig
+ 3.501000000e-07 V_hig
+ 3.501010000e-07 V_hig
+ 3.502000000e-07 V_hig
+ 3.502010000e-07 V_hig
+ 3.503000000e-07 V_hig
+ 3.503010000e-07 V_hig
+ 3.504000000e-07 V_hig
+ 3.504010000e-07 V_hig
+ 3.505000000e-07 V_hig
+ 3.505010000e-07 V_hig
+ 3.506000000e-07 V_hig
+ 3.506010000e-07 V_hig
+ 3.507000000e-07 V_hig
+ 3.507010000e-07 V_hig
+ 3.508000000e-07 V_hig
+ 3.508010000e-07 V_hig
+ 3.509000000e-07 V_hig
+ 3.509010000e-07 V_low
+ 3.510000000e-07 V_low
+ 3.510010000e-07 V_low
+ 3.511000000e-07 V_low
+ 3.511010000e-07 V_low
+ 3.512000000e-07 V_low
+ 3.512010000e-07 V_low
+ 3.513000000e-07 V_low
+ 3.513010000e-07 V_low
+ 3.514000000e-07 V_low
+ 3.514010000e-07 V_low
+ 3.515000000e-07 V_low
+ 3.515010000e-07 V_low
+ 3.516000000e-07 V_low
+ 3.516010000e-07 V_low
+ 3.517000000e-07 V_low
+ 3.517010000e-07 V_low
+ 3.518000000e-07 V_low
+ 3.518010000e-07 V_low
+ 3.519000000e-07 V_low
+ 3.519010000e-07 V_hig
+ 3.520000000e-07 V_hig
+ 3.520010000e-07 V_hig
+ 3.521000000e-07 V_hig
+ 3.521010000e-07 V_hig
+ 3.522000000e-07 V_hig
+ 3.522010000e-07 V_hig
+ 3.523000000e-07 V_hig
+ 3.523010000e-07 V_hig
+ 3.524000000e-07 V_hig
+ 3.524010000e-07 V_hig
+ 3.525000000e-07 V_hig
+ 3.525010000e-07 V_hig
+ 3.526000000e-07 V_hig
+ 3.526010000e-07 V_hig
+ 3.527000000e-07 V_hig
+ 3.527010000e-07 V_hig
+ 3.528000000e-07 V_hig
+ 3.528010000e-07 V_hig
+ 3.529000000e-07 V_hig
+ 3.529010000e-07 V_hig
+ 3.530000000e-07 V_hig
+ 3.530010000e-07 V_hig
+ 3.531000000e-07 V_hig
+ 3.531010000e-07 V_hig
+ 3.532000000e-07 V_hig
+ 3.532010000e-07 V_hig
+ 3.533000000e-07 V_hig
+ 3.533010000e-07 V_hig
+ 3.534000000e-07 V_hig
+ 3.534010000e-07 V_hig
+ 3.535000000e-07 V_hig
+ 3.535010000e-07 V_hig
+ 3.536000000e-07 V_hig
+ 3.536010000e-07 V_hig
+ 3.537000000e-07 V_hig
+ 3.537010000e-07 V_hig
+ 3.538000000e-07 V_hig
+ 3.538010000e-07 V_hig
+ 3.539000000e-07 V_hig
+ 3.539010000e-07 V_hig
+ 3.540000000e-07 V_hig
+ 3.540010000e-07 V_hig
+ 3.541000000e-07 V_hig
+ 3.541010000e-07 V_hig
+ 3.542000000e-07 V_hig
+ 3.542010000e-07 V_hig
+ 3.543000000e-07 V_hig
+ 3.543010000e-07 V_hig
+ 3.544000000e-07 V_hig
+ 3.544010000e-07 V_hig
+ 3.545000000e-07 V_hig
+ 3.545010000e-07 V_hig
+ 3.546000000e-07 V_hig
+ 3.546010000e-07 V_hig
+ 3.547000000e-07 V_hig
+ 3.547010000e-07 V_hig
+ 3.548000000e-07 V_hig
+ 3.548010000e-07 V_hig
+ 3.549000000e-07 V_hig
+ 3.549010000e-07 V_low
+ 3.550000000e-07 V_low
+ 3.550010000e-07 V_low
+ 3.551000000e-07 V_low
+ 3.551010000e-07 V_low
+ 3.552000000e-07 V_low
+ 3.552010000e-07 V_low
+ 3.553000000e-07 V_low
+ 3.553010000e-07 V_low
+ 3.554000000e-07 V_low
+ 3.554010000e-07 V_low
+ 3.555000000e-07 V_low
+ 3.555010000e-07 V_low
+ 3.556000000e-07 V_low
+ 3.556010000e-07 V_low
+ 3.557000000e-07 V_low
+ 3.557010000e-07 V_low
+ 3.558000000e-07 V_low
+ 3.558010000e-07 V_low
+ 3.559000000e-07 V_low
+ 3.559010000e-07 V_low
+ 3.560000000e-07 V_low
+ 3.560010000e-07 V_low
+ 3.561000000e-07 V_low
+ 3.561010000e-07 V_low
+ 3.562000000e-07 V_low
+ 3.562010000e-07 V_low
+ 3.563000000e-07 V_low
+ 3.563010000e-07 V_low
+ 3.564000000e-07 V_low
+ 3.564010000e-07 V_low
+ 3.565000000e-07 V_low
+ 3.565010000e-07 V_low
+ 3.566000000e-07 V_low
+ 3.566010000e-07 V_low
+ 3.567000000e-07 V_low
+ 3.567010000e-07 V_low
+ 3.568000000e-07 V_low
+ 3.568010000e-07 V_low
+ 3.569000000e-07 V_low
+ 3.569010000e-07 V_low
+ 3.570000000e-07 V_low
+ 3.570010000e-07 V_low
+ 3.571000000e-07 V_low
+ 3.571010000e-07 V_low
+ 3.572000000e-07 V_low
+ 3.572010000e-07 V_low
+ 3.573000000e-07 V_low
+ 3.573010000e-07 V_low
+ 3.574000000e-07 V_low
+ 3.574010000e-07 V_low
+ 3.575000000e-07 V_low
+ 3.575010000e-07 V_low
+ 3.576000000e-07 V_low
+ 3.576010000e-07 V_low
+ 3.577000000e-07 V_low
+ 3.577010000e-07 V_low
+ 3.578000000e-07 V_low
+ 3.578010000e-07 V_low
+ 3.579000000e-07 V_low
+ 3.579010000e-07 V_hig
+ 3.580000000e-07 V_hig
+ 3.580010000e-07 V_hig
+ 3.581000000e-07 V_hig
+ 3.581010000e-07 V_hig
+ 3.582000000e-07 V_hig
+ 3.582010000e-07 V_hig
+ 3.583000000e-07 V_hig
+ 3.583010000e-07 V_hig
+ 3.584000000e-07 V_hig
+ 3.584010000e-07 V_hig
+ 3.585000000e-07 V_hig
+ 3.585010000e-07 V_hig
+ 3.586000000e-07 V_hig
+ 3.586010000e-07 V_hig
+ 3.587000000e-07 V_hig
+ 3.587010000e-07 V_hig
+ 3.588000000e-07 V_hig
+ 3.588010000e-07 V_hig
+ 3.589000000e-07 V_hig
+ 3.589010000e-07 V_hig
+ 3.590000000e-07 V_hig
+ 3.590010000e-07 V_hig
+ 3.591000000e-07 V_hig
+ 3.591010000e-07 V_hig
+ 3.592000000e-07 V_hig
+ 3.592010000e-07 V_hig
+ 3.593000000e-07 V_hig
+ 3.593010000e-07 V_hig
+ 3.594000000e-07 V_hig
+ 3.594010000e-07 V_hig
+ 3.595000000e-07 V_hig
+ 3.595010000e-07 V_hig
+ 3.596000000e-07 V_hig
+ 3.596010000e-07 V_hig
+ 3.597000000e-07 V_hig
+ 3.597010000e-07 V_hig
+ 3.598000000e-07 V_hig
+ 3.598010000e-07 V_hig
+ 3.599000000e-07 V_hig
+ 3.599010000e-07 V_hig
+ 3.600000000e-07 V_hig
+ 3.600010000e-07 V_hig
+ 3.601000000e-07 V_hig
+ 3.601010000e-07 V_hig
+ 3.602000000e-07 V_hig
+ 3.602010000e-07 V_hig
+ 3.603000000e-07 V_hig
+ 3.603010000e-07 V_hig
+ 3.604000000e-07 V_hig
+ 3.604010000e-07 V_hig
+ 3.605000000e-07 V_hig
+ 3.605010000e-07 V_hig
+ 3.606000000e-07 V_hig
+ 3.606010000e-07 V_hig
+ 3.607000000e-07 V_hig
+ 3.607010000e-07 V_hig
+ 3.608000000e-07 V_hig
+ 3.608010000e-07 V_hig
+ 3.609000000e-07 V_hig
+ 3.609010000e-07 V_hig
+ 3.610000000e-07 V_hig
+ 3.610010000e-07 V_hig
+ 3.611000000e-07 V_hig
+ 3.611010000e-07 V_hig
+ 3.612000000e-07 V_hig
+ 3.612010000e-07 V_hig
+ 3.613000000e-07 V_hig
+ 3.613010000e-07 V_hig
+ 3.614000000e-07 V_hig
+ 3.614010000e-07 V_hig
+ 3.615000000e-07 V_hig
+ 3.615010000e-07 V_hig
+ 3.616000000e-07 V_hig
+ 3.616010000e-07 V_hig
+ 3.617000000e-07 V_hig
+ 3.617010000e-07 V_hig
+ 3.618000000e-07 V_hig
+ 3.618010000e-07 V_hig
+ 3.619000000e-07 V_hig
+ 3.619010000e-07 V_low
+ 3.620000000e-07 V_low
+ 3.620010000e-07 V_low
+ 3.621000000e-07 V_low
+ 3.621010000e-07 V_low
+ 3.622000000e-07 V_low
+ 3.622010000e-07 V_low
+ 3.623000000e-07 V_low
+ 3.623010000e-07 V_low
+ 3.624000000e-07 V_low
+ 3.624010000e-07 V_low
+ 3.625000000e-07 V_low
+ 3.625010000e-07 V_low
+ 3.626000000e-07 V_low
+ 3.626010000e-07 V_low
+ 3.627000000e-07 V_low
+ 3.627010000e-07 V_low
+ 3.628000000e-07 V_low
+ 3.628010000e-07 V_low
+ 3.629000000e-07 V_low
+ 3.629010000e-07 V_low
+ 3.630000000e-07 V_low
+ 3.630010000e-07 V_low
+ 3.631000000e-07 V_low
+ 3.631010000e-07 V_low
+ 3.632000000e-07 V_low
+ 3.632010000e-07 V_low
+ 3.633000000e-07 V_low
+ 3.633010000e-07 V_low
+ 3.634000000e-07 V_low
+ 3.634010000e-07 V_low
+ 3.635000000e-07 V_low
+ 3.635010000e-07 V_low
+ 3.636000000e-07 V_low
+ 3.636010000e-07 V_low
+ 3.637000000e-07 V_low
+ 3.637010000e-07 V_low
+ 3.638000000e-07 V_low
+ 3.638010000e-07 V_low
+ 3.639000000e-07 V_low
+ 3.639010000e-07 V_low
+ 3.640000000e-07 V_low
+ 3.640010000e-07 V_low
+ 3.641000000e-07 V_low
+ 3.641010000e-07 V_low
+ 3.642000000e-07 V_low
+ 3.642010000e-07 V_low
+ 3.643000000e-07 V_low
+ 3.643010000e-07 V_low
+ 3.644000000e-07 V_low
+ 3.644010000e-07 V_low
+ 3.645000000e-07 V_low
+ 3.645010000e-07 V_low
+ 3.646000000e-07 V_low
+ 3.646010000e-07 V_low
+ 3.647000000e-07 V_low
+ 3.647010000e-07 V_low
+ 3.648000000e-07 V_low
+ 3.648010000e-07 V_low
+ 3.649000000e-07 V_low
+ 3.649010000e-07 V_hig
+ 3.650000000e-07 V_hig
+ 3.650010000e-07 V_hig
+ 3.651000000e-07 V_hig
+ 3.651010000e-07 V_hig
+ 3.652000000e-07 V_hig
+ 3.652010000e-07 V_hig
+ 3.653000000e-07 V_hig
+ 3.653010000e-07 V_hig
+ 3.654000000e-07 V_hig
+ 3.654010000e-07 V_hig
+ 3.655000000e-07 V_hig
+ 3.655010000e-07 V_hig
+ 3.656000000e-07 V_hig
+ 3.656010000e-07 V_hig
+ 3.657000000e-07 V_hig
+ 3.657010000e-07 V_hig
+ 3.658000000e-07 V_hig
+ 3.658010000e-07 V_hig
+ 3.659000000e-07 V_hig
+ 3.659010000e-07 V_hig
+ 3.660000000e-07 V_hig
+ 3.660010000e-07 V_hig
+ 3.661000000e-07 V_hig
+ 3.661010000e-07 V_hig
+ 3.662000000e-07 V_hig
+ 3.662010000e-07 V_hig
+ 3.663000000e-07 V_hig
+ 3.663010000e-07 V_hig
+ 3.664000000e-07 V_hig
+ 3.664010000e-07 V_hig
+ 3.665000000e-07 V_hig
+ 3.665010000e-07 V_hig
+ 3.666000000e-07 V_hig
+ 3.666010000e-07 V_hig
+ 3.667000000e-07 V_hig
+ 3.667010000e-07 V_hig
+ 3.668000000e-07 V_hig
+ 3.668010000e-07 V_hig
+ 3.669000000e-07 V_hig
+ 3.669010000e-07 V_hig
+ 3.670000000e-07 V_hig
+ 3.670010000e-07 V_hig
+ 3.671000000e-07 V_hig
+ 3.671010000e-07 V_hig
+ 3.672000000e-07 V_hig
+ 3.672010000e-07 V_hig
+ 3.673000000e-07 V_hig
+ 3.673010000e-07 V_hig
+ 3.674000000e-07 V_hig
+ 3.674010000e-07 V_hig
+ 3.675000000e-07 V_hig
+ 3.675010000e-07 V_hig
+ 3.676000000e-07 V_hig
+ 3.676010000e-07 V_hig
+ 3.677000000e-07 V_hig
+ 3.677010000e-07 V_hig
+ 3.678000000e-07 V_hig
+ 3.678010000e-07 V_hig
+ 3.679000000e-07 V_hig
+ 3.679010000e-07 V_hig
+ 3.680000000e-07 V_hig
+ 3.680010000e-07 V_hig
+ 3.681000000e-07 V_hig
+ 3.681010000e-07 V_hig
+ 3.682000000e-07 V_hig
+ 3.682010000e-07 V_hig
+ 3.683000000e-07 V_hig
+ 3.683010000e-07 V_hig
+ 3.684000000e-07 V_hig
+ 3.684010000e-07 V_hig
+ 3.685000000e-07 V_hig
+ 3.685010000e-07 V_hig
+ 3.686000000e-07 V_hig
+ 3.686010000e-07 V_hig
+ 3.687000000e-07 V_hig
+ 3.687010000e-07 V_hig
+ 3.688000000e-07 V_hig
+ 3.688010000e-07 V_hig
+ 3.689000000e-07 V_hig
+ 3.689010000e-07 V_low
+ 3.690000000e-07 V_low
+ 3.690010000e-07 V_low
+ 3.691000000e-07 V_low
+ 3.691010000e-07 V_low
+ 3.692000000e-07 V_low
+ 3.692010000e-07 V_low
+ 3.693000000e-07 V_low
+ 3.693010000e-07 V_low
+ 3.694000000e-07 V_low
+ 3.694010000e-07 V_low
+ 3.695000000e-07 V_low
+ 3.695010000e-07 V_low
+ 3.696000000e-07 V_low
+ 3.696010000e-07 V_low
+ 3.697000000e-07 V_low
+ 3.697010000e-07 V_low
+ 3.698000000e-07 V_low
+ 3.698010000e-07 V_low
+ 3.699000000e-07 V_low
+ 3.699010000e-07 V_hig
+ 3.700000000e-07 V_hig
+ 3.700010000e-07 V_hig
+ 3.701000000e-07 V_hig
+ 3.701010000e-07 V_hig
+ 3.702000000e-07 V_hig
+ 3.702010000e-07 V_hig
+ 3.703000000e-07 V_hig
+ 3.703010000e-07 V_hig
+ 3.704000000e-07 V_hig
+ 3.704010000e-07 V_hig
+ 3.705000000e-07 V_hig
+ 3.705010000e-07 V_hig
+ 3.706000000e-07 V_hig
+ 3.706010000e-07 V_hig
+ 3.707000000e-07 V_hig
+ 3.707010000e-07 V_hig
+ 3.708000000e-07 V_hig
+ 3.708010000e-07 V_hig
+ 3.709000000e-07 V_hig
+ 3.709010000e-07 V_hig
+ 3.710000000e-07 V_hig
+ 3.710010000e-07 V_hig
+ 3.711000000e-07 V_hig
+ 3.711010000e-07 V_hig
+ 3.712000000e-07 V_hig
+ 3.712010000e-07 V_hig
+ 3.713000000e-07 V_hig
+ 3.713010000e-07 V_hig
+ 3.714000000e-07 V_hig
+ 3.714010000e-07 V_hig
+ 3.715000000e-07 V_hig
+ 3.715010000e-07 V_hig
+ 3.716000000e-07 V_hig
+ 3.716010000e-07 V_hig
+ 3.717000000e-07 V_hig
+ 3.717010000e-07 V_hig
+ 3.718000000e-07 V_hig
+ 3.718010000e-07 V_hig
+ 3.719000000e-07 V_hig
+ 3.719010000e-07 V_hig
+ 3.720000000e-07 V_hig
+ 3.720010000e-07 V_hig
+ 3.721000000e-07 V_hig
+ 3.721010000e-07 V_hig
+ 3.722000000e-07 V_hig
+ 3.722010000e-07 V_hig
+ 3.723000000e-07 V_hig
+ 3.723010000e-07 V_hig
+ 3.724000000e-07 V_hig
+ 3.724010000e-07 V_hig
+ 3.725000000e-07 V_hig
+ 3.725010000e-07 V_hig
+ 3.726000000e-07 V_hig
+ 3.726010000e-07 V_hig
+ 3.727000000e-07 V_hig
+ 3.727010000e-07 V_hig
+ 3.728000000e-07 V_hig
+ 3.728010000e-07 V_hig
+ 3.729000000e-07 V_hig
+ 3.729010000e-07 V_hig
+ 3.730000000e-07 V_hig
+ 3.730010000e-07 V_hig
+ 3.731000000e-07 V_hig
+ 3.731010000e-07 V_hig
+ 3.732000000e-07 V_hig
+ 3.732010000e-07 V_hig
+ 3.733000000e-07 V_hig
+ 3.733010000e-07 V_hig
+ 3.734000000e-07 V_hig
+ 3.734010000e-07 V_hig
+ 3.735000000e-07 V_hig
+ 3.735010000e-07 V_hig
+ 3.736000000e-07 V_hig
+ 3.736010000e-07 V_hig
+ 3.737000000e-07 V_hig
+ 3.737010000e-07 V_hig
+ 3.738000000e-07 V_hig
+ 3.738010000e-07 V_hig
+ 3.739000000e-07 V_hig
+ 3.739010000e-07 V_hig
+ 3.740000000e-07 V_hig
+ 3.740010000e-07 V_hig
+ 3.741000000e-07 V_hig
+ 3.741010000e-07 V_hig
+ 3.742000000e-07 V_hig
+ 3.742010000e-07 V_hig
+ 3.743000000e-07 V_hig
+ 3.743010000e-07 V_hig
+ 3.744000000e-07 V_hig
+ 3.744010000e-07 V_hig
+ 3.745000000e-07 V_hig
+ 3.745010000e-07 V_hig
+ 3.746000000e-07 V_hig
+ 3.746010000e-07 V_hig
+ 3.747000000e-07 V_hig
+ 3.747010000e-07 V_hig
+ 3.748000000e-07 V_hig
+ 3.748010000e-07 V_hig
+ 3.749000000e-07 V_hig
+ 3.749010000e-07 V_hig
+ 3.750000000e-07 V_hig
+ 3.750010000e-07 V_hig
+ 3.751000000e-07 V_hig
+ 3.751010000e-07 V_hig
+ 3.752000000e-07 V_hig
+ 3.752010000e-07 V_hig
+ 3.753000000e-07 V_hig
+ 3.753010000e-07 V_hig
+ 3.754000000e-07 V_hig
+ 3.754010000e-07 V_hig
+ 3.755000000e-07 V_hig
+ 3.755010000e-07 V_hig
+ 3.756000000e-07 V_hig
+ 3.756010000e-07 V_hig
+ 3.757000000e-07 V_hig
+ 3.757010000e-07 V_hig
+ 3.758000000e-07 V_hig
+ 3.758010000e-07 V_hig
+ 3.759000000e-07 V_hig
+ 3.759010000e-07 V_hig
+ 3.760000000e-07 V_hig
+ 3.760010000e-07 V_hig
+ 3.761000000e-07 V_hig
+ 3.761010000e-07 V_hig
+ 3.762000000e-07 V_hig
+ 3.762010000e-07 V_hig
+ 3.763000000e-07 V_hig
+ 3.763010000e-07 V_hig
+ 3.764000000e-07 V_hig
+ 3.764010000e-07 V_hig
+ 3.765000000e-07 V_hig
+ 3.765010000e-07 V_hig
+ 3.766000000e-07 V_hig
+ 3.766010000e-07 V_hig
+ 3.767000000e-07 V_hig
+ 3.767010000e-07 V_hig
+ 3.768000000e-07 V_hig
+ 3.768010000e-07 V_hig
+ 3.769000000e-07 V_hig
+ 3.769010000e-07 V_low
+ 3.770000000e-07 V_low
+ 3.770010000e-07 V_low
+ 3.771000000e-07 V_low
+ 3.771010000e-07 V_low
+ 3.772000000e-07 V_low
+ 3.772010000e-07 V_low
+ 3.773000000e-07 V_low
+ 3.773010000e-07 V_low
+ 3.774000000e-07 V_low
+ 3.774010000e-07 V_low
+ 3.775000000e-07 V_low
+ 3.775010000e-07 V_low
+ 3.776000000e-07 V_low
+ 3.776010000e-07 V_low
+ 3.777000000e-07 V_low
+ 3.777010000e-07 V_low
+ 3.778000000e-07 V_low
+ 3.778010000e-07 V_low
+ 3.779000000e-07 V_low
+ 3.779010000e-07 V_hig
+ 3.780000000e-07 V_hig
+ 3.780010000e-07 V_hig
+ 3.781000000e-07 V_hig
+ 3.781010000e-07 V_hig
+ 3.782000000e-07 V_hig
+ 3.782010000e-07 V_hig
+ 3.783000000e-07 V_hig
+ 3.783010000e-07 V_hig
+ 3.784000000e-07 V_hig
+ 3.784010000e-07 V_hig
+ 3.785000000e-07 V_hig
+ 3.785010000e-07 V_hig
+ 3.786000000e-07 V_hig
+ 3.786010000e-07 V_hig
+ 3.787000000e-07 V_hig
+ 3.787010000e-07 V_hig
+ 3.788000000e-07 V_hig
+ 3.788010000e-07 V_hig
+ 3.789000000e-07 V_hig
+ 3.789010000e-07 V_hig
+ 3.790000000e-07 V_hig
+ 3.790010000e-07 V_hig
+ 3.791000000e-07 V_hig
+ 3.791010000e-07 V_hig
+ 3.792000000e-07 V_hig
+ 3.792010000e-07 V_hig
+ 3.793000000e-07 V_hig
+ 3.793010000e-07 V_hig
+ 3.794000000e-07 V_hig
+ 3.794010000e-07 V_hig
+ 3.795000000e-07 V_hig
+ 3.795010000e-07 V_hig
+ 3.796000000e-07 V_hig
+ 3.796010000e-07 V_hig
+ 3.797000000e-07 V_hig
+ 3.797010000e-07 V_hig
+ 3.798000000e-07 V_hig
+ 3.798010000e-07 V_hig
+ 3.799000000e-07 V_hig
+ 3.799010000e-07 V_hig
+ 3.800000000e-07 V_hig
+ 3.800010000e-07 V_hig
+ 3.801000000e-07 V_hig
+ 3.801010000e-07 V_hig
+ 3.802000000e-07 V_hig
+ 3.802010000e-07 V_hig
+ 3.803000000e-07 V_hig
+ 3.803010000e-07 V_hig
+ 3.804000000e-07 V_hig
+ 3.804010000e-07 V_hig
+ 3.805000000e-07 V_hig
+ 3.805010000e-07 V_hig
+ 3.806000000e-07 V_hig
+ 3.806010000e-07 V_hig
+ 3.807000000e-07 V_hig
+ 3.807010000e-07 V_hig
+ 3.808000000e-07 V_hig
+ 3.808010000e-07 V_hig
+ 3.809000000e-07 V_hig
+ 3.809010000e-07 V_low
+ 3.810000000e-07 V_low
+ 3.810010000e-07 V_low
+ 3.811000000e-07 V_low
+ 3.811010000e-07 V_low
+ 3.812000000e-07 V_low
+ 3.812010000e-07 V_low
+ 3.813000000e-07 V_low
+ 3.813010000e-07 V_low
+ 3.814000000e-07 V_low
+ 3.814010000e-07 V_low
+ 3.815000000e-07 V_low
+ 3.815010000e-07 V_low
+ 3.816000000e-07 V_low
+ 3.816010000e-07 V_low
+ 3.817000000e-07 V_low
+ 3.817010000e-07 V_low
+ 3.818000000e-07 V_low
+ 3.818010000e-07 V_low
+ 3.819000000e-07 V_low
+ 3.819010000e-07 V_hig
+ 3.820000000e-07 V_hig
+ 3.820010000e-07 V_hig
+ 3.821000000e-07 V_hig
+ 3.821010000e-07 V_hig
+ 3.822000000e-07 V_hig
+ 3.822010000e-07 V_hig
+ 3.823000000e-07 V_hig
+ 3.823010000e-07 V_hig
+ 3.824000000e-07 V_hig
+ 3.824010000e-07 V_hig
+ 3.825000000e-07 V_hig
+ 3.825010000e-07 V_hig
+ 3.826000000e-07 V_hig
+ 3.826010000e-07 V_hig
+ 3.827000000e-07 V_hig
+ 3.827010000e-07 V_hig
+ 3.828000000e-07 V_hig
+ 3.828010000e-07 V_hig
+ 3.829000000e-07 V_hig
+ 3.829010000e-07 V_hig
+ 3.830000000e-07 V_hig
+ 3.830010000e-07 V_hig
+ 3.831000000e-07 V_hig
+ 3.831010000e-07 V_hig
+ 3.832000000e-07 V_hig
+ 3.832010000e-07 V_hig
+ 3.833000000e-07 V_hig
+ 3.833010000e-07 V_hig
+ 3.834000000e-07 V_hig
+ 3.834010000e-07 V_hig
+ 3.835000000e-07 V_hig
+ 3.835010000e-07 V_hig
+ 3.836000000e-07 V_hig
+ 3.836010000e-07 V_hig
+ 3.837000000e-07 V_hig
+ 3.837010000e-07 V_hig
+ 3.838000000e-07 V_hig
+ 3.838010000e-07 V_hig
+ 3.839000000e-07 V_hig
+ 3.839010000e-07 V_low
+ 3.840000000e-07 V_low
+ 3.840010000e-07 V_low
+ 3.841000000e-07 V_low
+ 3.841010000e-07 V_low
+ 3.842000000e-07 V_low
+ 3.842010000e-07 V_low
+ 3.843000000e-07 V_low
+ 3.843010000e-07 V_low
+ 3.844000000e-07 V_low
+ 3.844010000e-07 V_low
+ 3.845000000e-07 V_low
+ 3.845010000e-07 V_low
+ 3.846000000e-07 V_low
+ 3.846010000e-07 V_low
+ 3.847000000e-07 V_low
+ 3.847010000e-07 V_low
+ 3.848000000e-07 V_low
+ 3.848010000e-07 V_low
+ 3.849000000e-07 V_low
+ 3.849010000e-07 V_low
+ 3.850000000e-07 V_low
+ 3.850010000e-07 V_low
+ 3.851000000e-07 V_low
+ 3.851010000e-07 V_low
+ 3.852000000e-07 V_low
+ 3.852010000e-07 V_low
+ 3.853000000e-07 V_low
+ 3.853010000e-07 V_low
+ 3.854000000e-07 V_low
+ 3.854010000e-07 V_low
+ 3.855000000e-07 V_low
+ 3.855010000e-07 V_low
+ 3.856000000e-07 V_low
+ 3.856010000e-07 V_low
+ 3.857000000e-07 V_low
+ 3.857010000e-07 V_low
+ 3.858000000e-07 V_low
+ 3.858010000e-07 V_low
+ 3.859000000e-07 V_low
+ 3.859010000e-07 V_low
+ 3.860000000e-07 V_low
+ 3.860010000e-07 V_low
+ 3.861000000e-07 V_low
+ 3.861010000e-07 V_low
+ 3.862000000e-07 V_low
+ 3.862010000e-07 V_low
+ 3.863000000e-07 V_low
+ 3.863010000e-07 V_low
+ 3.864000000e-07 V_low
+ 3.864010000e-07 V_low
+ 3.865000000e-07 V_low
+ 3.865010000e-07 V_low
+ 3.866000000e-07 V_low
+ 3.866010000e-07 V_low
+ 3.867000000e-07 V_low
+ 3.867010000e-07 V_low
+ 3.868000000e-07 V_low
+ 3.868010000e-07 V_low
+ 3.869000000e-07 V_low
+ 3.869010000e-07 V_hig
+ 3.870000000e-07 V_hig
+ 3.870010000e-07 V_hig
+ 3.871000000e-07 V_hig
+ 3.871010000e-07 V_hig
+ 3.872000000e-07 V_hig
+ 3.872010000e-07 V_hig
+ 3.873000000e-07 V_hig
+ 3.873010000e-07 V_hig
+ 3.874000000e-07 V_hig
+ 3.874010000e-07 V_hig
+ 3.875000000e-07 V_hig
+ 3.875010000e-07 V_hig
+ 3.876000000e-07 V_hig
+ 3.876010000e-07 V_hig
+ 3.877000000e-07 V_hig
+ 3.877010000e-07 V_hig
+ 3.878000000e-07 V_hig
+ 3.878010000e-07 V_hig
+ 3.879000000e-07 V_hig
+ 3.879010000e-07 V_low
+ 3.880000000e-07 V_low
+ 3.880010000e-07 V_low
+ 3.881000000e-07 V_low
+ 3.881010000e-07 V_low
+ 3.882000000e-07 V_low
+ 3.882010000e-07 V_low
+ 3.883000000e-07 V_low
+ 3.883010000e-07 V_low
+ 3.884000000e-07 V_low
+ 3.884010000e-07 V_low
+ 3.885000000e-07 V_low
+ 3.885010000e-07 V_low
+ 3.886000000e-07 V_low
+ 3.886010000e-07 V_low
+ 3.887000000e-07 V_low
+ 3.887010000e-07 V_low
+ 3.888000000e-07 V_low
+ 3.888010000e-07 V_low
+ 3.889000000e-07 V_low
+ 3.889010000e-07 V_low
+ 3.890000000e-07 V_low
+ 3.890010000e-07 V_low
+ 3.891000000e-07 V_low
+ 3.891010000e-07 V_low
+ 3.892000000e-07 V_low
+ 3.892010000e-07 V_low
+ 3.893000000e-07 V_low
+ 3.893010000e-07 V_low
+ 3.894000000e-07 V_low
+ 3.894010000e-07 V_low
+ 3.895000000e-07 V_low
+ 3.895010000e-07 V_low
+ 3.896000000e-07 V_low
+ 3.896010000e-07 V_low
+ 3.897000000e-07 V_low
+ 3.897010000e-07 V_low
+ 3.898000000e-07 V_low
+ 3.898010000e-07 V_low
+ 3.899000000e-07 V_low
+ 3.899010000e-07 V_low
+ 3.900000000e-07 V_low
+ 3.900010000e-07 V_low
+ 3.901000000e-07 V_low
+ 3.901010000e-07 V_low
+ 3.902000000e-07 V_low
+ 3.902010000e-07 V_low
+ 3.903000000e-07 V_low
+ 3.903010000e-07 V_low
+ 3.904000000e-07 V_low
+ 3.904010000e-07 V_low
+ 3.905000000e-07 V_low
+ 3.905010000e-07 V_low
+ 3.906000000e-07 V_low
+ 3.906010000e-07 V_low
+ 3.907000000e-07 V_low
+ 3.907010000e-07 V_low
+ 3.908000000e-07 V_low
+ 3.908010000e-07 V_low
+ 3.909000000e-07 V_low
+ 3.909010000e-07 V_hig
+ 3.910000000e-07 V_hig
+ 3.910010000e-07 V_hig
+ 3.911000000e-07 V_hig
+ 3.911010000e-07 V_hig
+ 3.912000000e-07 V_hig
+ 3.912010000e-07 V_hig
+ 3.913000000e-07 V_hig
+ 3.913010000e-07 V_hig
+ 3.914000000e-07 V_hig
+ 3.914010000e-07 V_hig
+ 3.915000000e-07 V_hig
+ 3.915010000e-07 V_hig
+ 3.916000000e-07 V_hig
+ 3.916010000e-07 V_hig
+ 3.917000000e-07 V_hig
+ 3.917010000e-07 V_hig
+ 3.918000000e-07 V_hig
+ 3.918010000e-07 V_hig
+ 3.919000000e-07 V_hig
+ 3.919010000e-07 V_hig
+ 3.920000000e-07 V_hig
+ 3.920010000e-07 V_hig
+ 3.921000000e-07 V_hig
+ 3.921010000e-07 V_hig
+ 3.922000000e-07 V_hig
+ 3.922010000e-07 V_hig
+ 3.923000000e-07 V_hig
+ 3.923010000e-07 V_hig
+ 3.924000000e-07 V_hig
+ 3.924010000e-07 V_hig
+ 3.925000000e-07 V_hig
+ 3.925010000e-07 V_hig
+ 3.926000000e-07 V_hig
+ 3.926010000e-07 V_hig
+ 3.927000000e-07 V_hig
+ 3.927010000e-07 V_hig
+ 3.928000000e-07 V_hig
+ 3.928010000e-07 V_hig
+ 3.929000000e-07 V_hig
+ 3.929010000e-07 V_low
+ 3.930000000e-07 V_low
+ 3.930010000e-07 V_low
+ 3.931000000e-07 V_low
+ 3.931010000e-07 V_low
+ 3.932000000e-07 V_low
+ 3.932010000e-07 V_low
+ 3.933000000e-07 V_low
+ 3.933010000e-07 V_low
+ 3.934000000e-07 V_low
+ 3.934010000e-07 V_low
+ 3.935000000e-07 V_low
+ 3.935010000e-07 V_low
+ 3.936000000e-07 V_low
+ 3.936010000e-07 V_low
+ 3.937000000e-07 V_low
+ 3.937010000e-07 V_low
+ 3.938000000e-07 V_low
+ 3.938010000e-07 V_low
+ 3.939000000e-07 V_low
+ 3.939010000e-07 V_low
+ 3.940000000e-07 V_low
+ 3.940010000e-07 V_low
+ 3.941000000e-07 V_low
+ 3.941010000e-07 V_low
+ 3.942000000e-07 V_low
+ 3.942010000e-07 V_low
+ 3.943000000e-07 V_low
+ 3.943010000e-07 V_low
+ 3.944000000e-07 V_low
+ 3.944010000e-07 V_low
+ 3.945000000e-07 V_low
+ 3.945010000e-07 V_low
+ 3.946000000e-07 V_low
+ 3.946010000e-07 V_low
+ 3.947000000e-07 V_low
+ 3.947010000e-07 V_low
+ 3.948000000e-07 V_low
+ 3.948010000e-07 V_low
+ 3.949000000e-07 V_low
+ 3.949010000e-07 V_hig
+ 3.950000000e-07 V_hig
+ 3.950010000e-07 V_hig
+ 3.951000000e-07 V_hig
+ 3.951010000e-07 V_hig
+ 3.952000000e-07 V_hig
+ 3.952010000e-07 V_hig
+ 3.953000000e-07 V_hig
+ 3.953010000e-07 V_hig
+ 3.954000000e-07 V_hig
+ 3.954010000e-07 V_hig
+ 3.955000000e-07 V_hig
+ 3.955010000e-07 V_hig
+ 3.956000000e-07 V_hig
+ 3.956010000e-07 V_hig
+ 3.957000000e-07 V_hig
+ 3.957010000e-07 V_hig
+ 3.958000000e-07 V_hig
+ 3.958010000e-07 V_hig
+ 3.959000000e-07 V_hig
+ 3.959010000e-07 V_hig
+ 3.960000000e-07 V_hig
+ 3.960010000e-07 V_hig
+ 3.961000000e-07 V_hig
+ 3.961010000e-07 V_hig
+ 3.962000000e-07 V_hig
+ 3.962010000e-07 V_hig
+ 3.963000000e-07 V_hig
+ 3.963010000e-07 V_hig
+ 3.964000000e-07 V_hig
+ 3.964010000e-07 V_hig
+ 3.965000000e-07 V_hig
+ 3.965010000e-07 V_hig
+ 3.966000000e-07 V_hig
+ 3.966010000e-07 V_hig
+ 3.967000000e-07 V_hig
+ 3.967010000e-07 V_hig
+ 3.968000000e-07 V_hig
+ 3.968010000e-07 V_hig
+ 3.969000000e-07 V_hig
+ 3.969010000e-07 V_hig
+ 3.970000000e-07 V_hig
+ 3.970010000e-07 V_hig
+ 3.971000000e-07 V_hig
+ 3.971010000e-07 V_hig
+ 3.972000000e-07 V_hig
+ 3.972010000e-07 V_hig
+ 3.973000000e-07 V_hig
+ 3.973010000e-07 V_hig
+ 3.974000000e-07 V_hig
+ 3.974010000e-07 V_hig
+ 3.975000000e-07 V_hig
+ 3.975010000e-07 V_hig
+ 3.976000000e-07 V_hig
+ 3.976010000e-07 V_hig
+ 3.977000000e-07 V_hig
+ 3.977010000e-07 V_hig
+ 3.978000000e-07 V_hig
+ 3.978010000e-07 V_hig
+ 3.979000000e-07 V_hig
+ 3.979010000e-07 V_hig
+ 3.980000000e-07 V_hig
+ 3.980010000e-07 V_hig
+ 3.981000000e-07 V_hig
+ 3.981010000e-07 V_hig
+ 3.982000000e-07 V_hig
+ 3.982010000e-07 V_hig
+ 3.983000000e-07 V_hig
+ 3.983010000e-07 V_hig
+ 3.984000000e-07 V_hig
+ 3.984010000e-07 V_hig
+ 3.985000000e-07 V_hig
+ 3.985010000e-07 V_hig
+ 3.986000000e-07 V_hig
+ 3.986010000e-07 V_hig
+ 3.987000000e-07 V_hig
+ 3.987010000e-07 V_hig
+ 3.988000000e-07 V_hig
+ 3.988010000e-07 V_hig
+ 3.989000000e-07 V_hig
+ 3.989010000e-07 V_low
+ 3.990000000e-07 V_low
+ 3.990010000e-07 V_low
+ 3.991000000e-07 V_low
+ 3.991010000e-07 V_low
+ 3.992000000e-07 V_low
+ 3.992010000e-07 V_low
+ 3.993000000e-07 V_low
+ 3.993010000e-07 V_low
+ 3.994000000e-07 V_low
+ 3.994010000e-07 V_low
+ 3.995000000e-07 V_low
+ 3.995010000e-07 V_low
+ 3.996000000e-07 V_low
+ 3.996010000e-07 V_low
+ 3.997000000e-07 V_low
+ 3.997010000e-07 V_low
+ 3.998000000e-07 V_low
+ 3.998010000e-07 V_low
+ 3.999000000e-07 V_low
+ 3.999010000e-07 V_low
+ 4.000000000e-07 V_low
+ 4.000010000e-07 V_low
+ 4.001000000e-07 V_low
+ 4.001010000e-07 V_low
+ 4.002000000e-07 V_low
+ 4.002010000e-07 V_low
+ 4.003000000e-07 V_low
+ 4.003010000e-07 V_low
+ 4.004000000e-07 V_low
+ 4.004010000e-07 V_low
+ 4.005000000e-07 V_low
+ 4.005010000e-07 V_low
+ 4.006000000e-07 V_low
+ 4.006010000e-07 V_low
+ 4.007000000e-07 V_low
+ 4.007010000e-07 V_low
+ 4.008000000e-07 V_low
+ 4.008010000e-07 V_low
+ 4.009000000e-07 V_low
+ 4.009010000e-07 V_hig
+ 4.010000000e-07 V_hig
+ 4.010010000e-07 V_hig
+ 4.011000000e-07 V_hig
+ 4.011010000e-07 V_hig
+ 4.012000000e-07 V_hig
+ 4.012010000e-07 V_hig
+ 4.013000000e-07 V_hig
+ 4.013010000e-07 V_hig
+ 4.014000000e-07 V_hig
+ 4.014010000e-07 V_hig
+ 4.015000000e-07 V_hig
+ 4.015010000e-07 V_hig
+ 4.016000000e-07 V_hig
+ 4.016010000e-07 V_hig
+ 4.017000000e-07 V_hig
+ 4.017010000e-07 V_hig
+ 4.018000000e-07 V_hig
+ 4.018010000e-07 V_hig
+ 4.019000000e-07 V_hig
+ 4.019010000e-07 V_low
+ 4.020000000e-07 V_low
+ 4.020010000e-07 V_low
+ 4.021000000e-07 V_low
+ 4.021010000e-07 V_low
+ 4.022000000e-07 V_low
+ 4.022010000e-07 V_low
+ 4.023000000e-07 V_low
+ 4.023010000e-07 V_low
+ 4.024000000e-07 V_low
+ 4.024010000e-07 V_low
+ 4.025000000e-07 V_low
+ 4.025010000e-07 V_low
+ 4.026000000e-07 V_low
+ 4.026010000e-07 V_low
+ 4.027000000e-07 V_low
+ 4.027010000e-07 V_low
+ 4.028000000e-07 V_low
+ 4.028010000e-07 V_low
+ 4.029000000e-07 V_low
+ 4.029010000e-07 V_low
+ 4.030000000e-07 V_low
+ 4.030010000e-07 V_low
+ 4.031000000e-07 V_low
+ 4.031010000e-07 V_low
+ 4.032000000e-07 V_low
+ 4.032010000e-07 V_low
+ 4.033000000e-07 V_low
+ 4.033010000e-07 V_low
+ 4.034000000e-07 V_low
+ 4.034010000e-07 V_low
+ 4.035000000e-07 V_low
+ 4.035010000e-07 V_low
+ 4.036000000e-07 V_low
+ 4.036010000e-07 V_low
+ 4.037000000e-07 V_low
+ 4.037010000e-07 V_low
+ 4.038000000e-07 V_low
+ 4.038010000e-07 V_low
+ 4.039000000e-07 V_low
+ 4.039010000e-07 V_low
+ 4.040000000e-07 V_low
+ 4.040010000e-07 V_low
+ 4.041000000e-07 V_low
+ 4.041010000e-07 V_low
+ 4.042000000e-07 V_low
+ 4.042010000e-07 V_low
+ 4.043000000e-07 V_low
+ 4.043010000e-07 V_low
+ 4.044000000e-07 V_low
+ 4.044010000e-07 V_low
+ 4.045000000e-07 V_low
+ 4.045010000e-07 V_low
+ 4.046000000e-07 V_low
+ 4.046010000e-07 V_low
+ 4.047000000e-07 V_low
+ 4.047010000e-07 V_low
+ 4.048000000e-07 V_low
+ 4.048010000e-07 V_low
+ 4.049000000e-07 V_low
+ 4.049010000e-07 V_hig
+ 4.050000000e-07 V_hig
+ 4.050010000e-07 V_hig
+ 4.051000000e-07 V_hig
+ 4.051010000e-07 V_hig
+ 4.052000000e-07 V_hig
+ 4.052010000e-07 V_hig
+ 4.053000000e-07 V_hig
+ 4.053010000e-07 V_hig
+ 4.054000000e-07 V_hig
+ 4.054010000e-07 V_hig
+ 4.055000000e-07 V_hig
+ 4.055010000e-07 V_hig
+ 4.056000000e-07 V_hig
+ 4.056010000e-07 V_hig
+ 4.057000000e-07 V_hig
+ 4.057010000e-07 V_hig
+ 4.058000000e-07 V_hig
+ 4.058010000e-07 V_hig
+ 4.059000000e-07 V_hig
+ 4.059010000e-07 V_low
+ 4.060000000e-07 V_low
+ 4.060010000e-07 V_low
+ 4.061000000e-07 V_low
+ 4.061010000e-07 V_low
+ 4.062000000e-07 V_low
+ 4.062010000e-07 V_low
+ 4.063000000e-07 V_low
+ 4.063010000e-07 V_low
+ 4.064000000e-07 V_low
+ 4.064010000e-07 V_low
+ 4.065000000e-07 V_low
+ 4.065010000e-07 V_low
+ 4.066000000e-07 V_low
+ 4.066010000e-07 V_low
+ 4.067000000e-07 V_low
+ 4.067010000e-07 V_low
+ 4.068000000e-07 V_low
+ 4.068010000e-07 V_low
+ 4.069000000e-07 V_low
+ 4.069010000e-07 V_hig
+ 4.070000000e-07 V_hig
+ 4.070010000e-07 V_hig
+ 4.071000000e-07 V_hig
+ 4.071010000e-07 V_hig
+ 4.072000000e-07 V_hig
+ 4.072010000e-07 V_hig
+ 4.073000000e-07 V_hig
+ 4.073010000e-07 V_hig
+ 4.074000000e-07 V_hig
+ 4.074010000e-07 V_hig
+ 4.075000000e-07 V_hig
+ 4.075010000e-07 V_hig
+ 4.076000000e-07 V_hig
+ 4.076010000e-07 V_hig
+ 4.077000000e-07 V_hig
+ 4.077010000e-07 V_hig
+ 4.078000000e-07 V_hig
+ 4.078010000e-07 V_hig
+ 4.079000000e-07 V_hig
+ 4.079010000e-07 V_low
+ 4.080000000e-07 V_low
+ 4.080010000e-07 V_low
+ 4.081000000e-07 V_low
+ 4.081010000e-07 V_low
+ 4.082000000e-07 V_low
+ 4.082010000e-07 V_low
+ 4.083000000e-07 V_low
+ 4.083010000e-07 V_low
+ 4.084000000e-07 V_low
+ 4.084010000e-07 V_low
+ 4.085000000e-07 V_low
+ 4.085010000e-07 V_low
+ 4.086000000e-07 V_low
+ 4.086010000e-07 V_low
+ 4.087000000e-07 V_low
+ 4.087010000e-07 V_low
+ 4.088000000e-07 V_low
+ 4.088010000e-07 V_low
+ 4.089000000e-07 V_low
+ 4.089010000e-07 V_low
+ 4.090000000e-07 V_low
+ 4.090010000e-07 V_low
+ 4.091000000e-07 V_low
+ 4.091010000e-07 V_low
+ 4.092000000e-07 V_low
+ 4.092010000e-07 V_low
+ 4.093000000e-07 V_low
+ 4.093010000e-07 V_low
+ 4.094000000e-07 V_low
+ 4.094010000e-07 V_low
+ 4.095000000e-07 V_low
+ 4.095010000e-07 V_low
+ 4.096000000e-07 V_low
+ 4.096010000e-07 V_low
+ 4.097000000e-07 V_low
+ 4.097010000e-07 V_low
+ 4.098000000e-07 V_low
+ 4.098010000e-07 V_low
+ 4.099000000e-07 V_low
+ 4.099010000e-07 V_hig
+ 4.100000000e-07 V_hig
+ 4.100010000e-07 V_hig
+ 4.101000000e-07 V_hig
+ 4.101010000e-07 V_hig
+ 4.102000000e-07 V_hig
+ 4.102010000e-07 V_hig
+ 4.103000000e-07 V_hig
+ 4.103010000e-07 V_hig
+ 4.104000000e-07 V_hig
+ 4.104010000e-07 V_hig
+ 4.105000000e-07 V_hig
+ 4.105010000e-07 V_hig
+ 4.106000000e-07 V_hig
+ 4.106010000e-07 V_hig
+ 4.107000000e-07 V_hig
+ 4.107010000e-07 V_hig
+ 4.108000000e-07 V_hig
+ 4.108010000e-07 V_hig
+ 4.109000000e-07 V_hig
+ 4.109010000e-07 V_low
+ 4.110000000e-07 V_low
+ 4.110010000e-07 V_low
+ 4.111000000e-07 V_low
+ 4.111010000e-07 V_low
+ 4.112000000e-07 V_low
+ 4.112010000e-07 V_low
+ 4.113000000e-07 V_low
+ 4.113010000e-07 V_low
+ 4.114000000e-07 V_low
+ 4.114010000e-07 V_low
+ 4.115000000e-07 V_low
+ 4.115010000e-07 V_low
+ 4.116000000e-07 V_low
+ 4.116010000e-07 V_low
+ 4.117000000e-07 V_low
+ 4.117010000e-07 V_low
+ 4.118000000e-07 V_low
+ 4.118010000e-07 V_low
+ 4.119000000e-07 V_low
+ 4.119010000e-07 V_low
+ 4.120000000e-07 V_low
+ 4.120010000e-07 V_low
+ 4.121000000e-07 V_low
+ 4.121010000e-07 V_low
+ 4.122000000e-07 V_low
+ 4.122010000e-07 V_low
+ 4.123000000e-07 V_low
+ 4.123010000e-07 V_low
+ 4.124000000e-07 V_low
+ 4.124010000e-07 V_low
+ 4.125000000e-07 V_low
+ 4.125010000e-07 V_low
+ 4.126000000e-07 V_low
+ 4.126010000e-07 V_low
+ 4.127000000e-07 V_low
+ 4.127010000e-07 V_low
+ 4.128000000e-07 V_low
+ 4.128010000e-07 V_low
+ 4.129000000e-07 V_low
+ 4.129010000e-07 V_low
+ 4.130000000e-07 V_low
+ 4.130010000e-07 V_low
+ 4.131000000e-07 V_low
+ 4.131010000e-07 V_low
+ 4.132000000e-07 V_low
+ 4.132010000e-07 V_low
+ 4.133000000e-07 V_low
+ 4.133010000e-07 V_low
+ 4.134000000e-07 V_low
+ 4.134010000e-07 V_low
+ 4.135000000e-07 V_low
+ 4.135010000e-07 V_low
+ 4.136000000e-07 V_low
+ 4.136010000e-07 V_low
+ 4.137000000e-07 V_low
+ 4.137010000e-07 V_low
+ 4.138000000e-07 V_low
+ 4.138010000e-07 V_low
+ 4.139000000e-07 V_low
+ 4.139010000e-07 V_hig
+ 4.140000000e-07 V_hig
+ 4.140010000e-07 V_hig
+ 4.141000000e-07 V_hig
+ 4.141010000e-07 V_hig
+ 4.142000000e-07 V_hig
+ 4.142010000e-07 V_hig
+ 4.143000000e-07 V_hig
+ 4.143010000e-07 V_hig
+ 4.144000000e-07 V_hig
+ 4.144010000e-07 V_hig
+ 4.145000000e-07 V_hig
+ 4.145010000e-07 V_hig
+ 4.146000000e-07 V_hig
+ 4.146010000e-07 V_hig
+ 4.147000000e-07 V_hig
+ 4.147010000e-07 V_hig
+ 4.148000000e-07 V_hig
+ 4.148010000e-07 V_hig
+ 4.149000000e-07 V_hig
+ 4.149010000e-07 V_hig
+ 4.150000000e-07 V_hig
+ 4.150010000e-07 V_hig
+ 4.151000000e-07 V_hig
+ 4.151010000e-07 V_hig
+ 4.152000000e-07 V_hig
+ 4.152010000e-07 V_hig
+ 4.153000000e-07 V_hig
+ 4.153010000e-07 V_hig
+ 4.154000000e-07 V_hig
+ 4.154010000e-07 V_hig
+ 4.155000000e-07 V_hig
+ 4.155010000e-07 V_hig
+ 4.156000000e-07 V_hig
+ 4.156010000e-07 V_hig
+ 4.157000000e-07 V_hig
+ 4.157010000e-07 V_hig
+ 4.158000000e-07 V_hig
+ 4.158010000e-07 V_hig
+ 4.159000000e-07 V_hig
+ 4.159010000e-07 V_hig
+ 4.160000000e-07 V_hig
+ 4.160010000e-07 V_hig
+ 4.161000000e-07 V_hig
+ 4.161010000e-07 V_hig
+ 4.162000000e-07 V_hig
+ 4.162010000e-07 V_hig
+ 4.163000000e-07 V_hig
+ 4.163010000e-07 V_hig
+ 4.164000000e-07 V_hig
+ 4.164010000e-07 V_hig
+ 4.165000000e-07 V_hig
+ 4.165010000e-07 V_hig
+ 4.166000000e-07 V_hig
+ 4.166010000e-07 V_hig
+ 4.167000000e-07 V_hig
+ 4.167010000e-07 V_hig
+ 4.168000000e-07 V_hig
+ 4.168010000e-07 V_hig
+ 4.169000000e-07 V_hig
+ 4.169010000e-07 V_low
+ 4.170000000e-07 V_low
+ 4.170010000e-07 V_low
+ 4.171000000e-07 V_low
+ 4.171010000e-07 V_low
+ 4.172000000e-07 V_low
+ 4.172010000e-07 V_low
+ 4.173000000e-07 V_low
+ 4.173010000e-07 V_low
+ 4.174000000e-07 V_low
+ 4.174010000e-07 V_low
+ 4.175000000e-07 V_low
+ 4.175010000e-07 V_low
+ 4.176000000e-07 V_low
+ 4.176010000e-07 V_low
+ 4.177000000e-07 V_low
+ 4.177010000e-07 V_low
+ 4.178000000e-07 V_low
+ 4.178010000e-07 V_low
+ 4.179000000e-07 V_low
+ 4.179010000e-07 V_low
+ 4.180000000e-07 V_low
+ 4.180010000e-07 V_low
+ 4.181000000e-07 V_low
+ 4.181010000e-07 V_low
+ 4.182000000e-07 V_low
+ 4.182010000e-07 V_low
+ 4.183000000e-07 V_low
+ 4.183010000e-07 V_low
+ 4.184000000e-07 V_low
+ 4.184010000e-07 V_low
+ 4.185000000e-07 V_low
+ 4.185010000e-07 V_low
+ 4.186000000e-07 V_low
+ 4.186010000e-07 V_low
+ 4.187000000e-07 V_low
+ 4.187010000e-07 V_low
+ 4.188000000e-07 V_low
+ 4.188010000e-07 V_low
+ 4.189000000e-07 V_low
+ 4.189010000e-07 V_hig
+ 4.190000000e-07 V_hig
+ 4.190010000e-07 V_hig
+ 4.191000000e-07 V_hig
+ 4.191010000e-07 V_hig
+ 4.192000000e-07 V_hig
+ 4.192010000e-07 V_hig
+ 4.193000000e-07 V_hig
+ 4.193010000e-07 V_hig
+ 4.194000000e-07 V_hig
+ 4.194010000e-07 V_hig
+ 4.195000000e-07 V_hig
+ 4.195010000e-07 V_hig
+ 4.196000000e-07 V_hig
+ 4.196010000e-07 V_hig
+ 4.197000000e-07 V_hig
+ 4.197010000e-07 V_hig
+ 4.198000000e-07 V_hig
+ 4.198010000e-07 V_hig
+ 4.199000000e-07 V_hig
+ 4.199010000e-07 V_hig
+ 4.200000000e-07 V_hig
+ 4.200010000e-07 V_hig
+ 4.201000000e-07 V_hig
+ 4.201010000e-07 V_hig
+ 4.202000000e-07 V_hig
+ 4.202010000e-07 V_hig
+ 4.203000000e-07 V_hig
+ 4.203010000e-07 V_hig
+ 4.204000000e-07 V_hig
+ 4.204010000e-07 V_hig
+ 4.205000000e-07 V_hig
+ 4.205010000e-07 V_hig
+ 4.206000000e-07 V_hig
+ 4.206010000e-07 V_hig
+ 4.207000000e-07 V_hig
+ 4.207010000e-07 V_hig
+ 4.208000000e-07 V_hig
+ 4.208010000e-07 V_hig
+ 4.209000000e-07 V_hig
+ 4.209010000e-07 V_low
+ 4.210000000e-07 V_low
+ 4.210010000e-07 V_low
+ 4.211000000e-07 V_low
+ 4.211010000e-07 V_low
+ 4.212000000e-07 V_low
+ 4.212010000e-07 V_low
+ 4.213000000e-07 V_low
+ 4.213010000e-07 V_low
+ 4.214000000e-07 V_low
+ 4.214010000e-07 V_low
+ 4.215000000e-07 V_low
+ 4.215010000e-07 V_low
+ 4.216000000e-07 V_low
+ 4.216010000e-07 V_low
+ 4.217000000e-07 V_low
+ 4.217010000e-07 V_low
+ 4.218000000e-07 V_low
+ 4.218010000e-07 V_low
+ 4.219000000e-07 V_low
+ 4.219010000e-07 V_low
+ 4.220000000e-07 V_low
+ 4.220010000e-07 V_low
+ 4.221000000e-07 V_low
+ 4.221010000e-07 V_low
+ 4.222000000e-07 V_low
+ 4.222010000e-07 V_low
+ 4.223000000e-07 V_low
+ 4.223010000e-07 V_low
+ 4.224000000e-07 V_low
+ 4.224010000e-07 V_low
+ 4.225000000e-07 V_low
+ 4.225010000e-07 V_low
+ 4.226000000e-07 V_low
+ 4.226010000e-07 V_low
+ 4.227000000e-07 V_low
+ 4.227010000e-07 V_low
+ 4.228000000e-07 V_low
+ 4.228010000e-07 V_low
+ 4.229000000e-07 V_low
+ 4.229010000e-07 V_low
+ 4.230000000e-07 V_low
+ 4.230010000e-07 V_low
+ 4.231000000e-07 V_low
+ 4.231010000e-07 V_low
+ 4.232000000e-07 V_low
+ 4.232010000e-07 V_low
+ 4.233000000e-07 V_low
+ 4.233010000e-07 V_low
+ 4.234000000e-07 V_low
+ 4.234010000e-07 V_low
+ 4.235000000e-07 V_low
+ 4.235010000e-07 V_low
+ 4.236000000e-07 V_low
+ 4.236010000e-07 V_low
+ 4.237000000e-07 V_low
+ 4.237010000e-07 V_low
+ 4.238000000e-07 V_low
+ 4.238010000e-07 V_low
+ 4.239000000e-07 V_low
+ 4.239010000e-07 V_hig
+ 4.240000000e-07 V_hig
+ 4.240010000e-07 V_hig
+ 4.241000000e-07 V_hig
+ 4.241010000e-07 V_hig
+ 4.242000000e-07 V_hig
+ 4.242010000e-07 V_hig
+ 4.243000000e-07 V_hig
+ 4.243010000e-07 V_hig
+ 4.244000000e-07 V_hig
+ 4.244010000e-07 V_hig
+ 4.245000000e-07 V_hig
+ 4.245010000e-07 V_hig
+ 4.246000000e-07 V_hig
+ 4.246010000e-07 V_hig
+ 4.247000000e-07 V_hig
+ 4.247010000e-07 V_hig
+ 4.248000000e-07 V_hig
+ 4.248010000e-07 V_hig
+ 4.249000000e-07 V_hig
+ 4.249010000e-07 V_low
+ 4.250000000e-07 V_low
+ 4.250010000e-07 V_low
+ 4.251000000e-07 V_low
+ 4.251010000e-07 V_low
+ 4.252000000e-07 V_low
+ 4.252010000e-07 V_low
+ 4.253000000e-07 V_low
+ 4.253010000e-07 V_low
+ 4.254000000e-07 V_low
+ 4.254010000e-07 V_low
+ 4.255000000e-07 V_low
+ 4.255010000e-07 V_low
+ 4.256000000e-07 V_low
+ 4.256010000e-07 V_low
+ 4.257000000e-07 V_low
+ 4.257010000e-07 V_low
+ 4.258000000e-07 V_low
+ 4.258010000e-07 V_low
+ 4.259000000e-07 V_low
+ 4.259010000e-07 V_hig
+ 4.260000000e-07 V_hig
+ 4.260010000e-07 V_hig
+ 4.261000000e-07 V_hig
+ 4.261010000e-07 V_hig
+ 4.262000000e-07 V_hig
+ 4.262010000e-07 V_hig
+ 4.263000000e-07 V_hig
+ 4.263010000e-07 V_hig
+ 4.264000000e-07 V_hig
+ 4.264010000e-07 V_hig
+ 4.265000000e-07 V_hig
+ 4.265010000e-07 V_hig
+ 4.266000000e-07 V_hig
+ 4.266010000e-07 V_hig
+ 4.267000000e-07 V_hig
+ 4.267010000e-07 V_hig
+ 4.268000000e-07 V_hig
+ 4.268010000e-07 V_hig
+ 4.269000000e-07 V_hig
+ 4.269010000e-07 V_hig
+ 4.270000000e-07 V_hig
+ 4.270010000e-07 V_hig
+ 4.271000000e-07 V_hig
+ 4.271010000e-07 V_hig
+ 4.272000000e-07 V_hig
+ 4.272010000e-07 V_hig
+ 4.273000000e-07 V_hig
+ 4.273010000e-07 V_hig
+ 4.274000000e-07 V_hig
+ 4.274010000e-07 V_hig
+ 4.275000000e-07 V_hig
+ 4.275010000e-07 V_hig
+ 4.276000000e-07 V_hig
+ 4.276010000e-07 V_hig
+ 4.277000000e-07 V_hig
+ 4.277010000e-07 V_hig
+ 4.278000000e-07 V_hig
+ 4.278010000e-07 V_hig
+ 4.279000000e-07 V_hig
+ 4.279010000e-07 V_hig
+ 4.280000000e-07 V_hig
+ 4.280010000e-07 V_hig
+ 4.281000000e-07 V_hig
+ 4.281010000e-07 V_hig
+ 4.282000000e-07 V_hig
+ 4.282010000e-07 V_hig
+ 4.283000000e-07 V_hig
+ 4.283010000e-07 V_hig
+ 4.284000000e-07 V_hig
+ 4.284010000e-07 V_hig
+ 4.285000000e-07 V_hig
+ 4.285010000e-07 V_hig
+ 4.286000000e-07 V_hig
+ 4.286010000e-07 V_hig
+ 4.287000000e-07 V_hig
+ 4.287010000e-07 V_hig
+ 4.288000000e-07 V_hig
+ 4.288010000e-07 V_hig
+ 4.289000000e-07 V_hig
+ 4.289010000e-07 V_hig
+ 4.290000000e-07 V_hig
+ 4.290010000e-07 V_hig
+ 4.291000000e-07 V_hig
+ 4.291010000e-07 V_hig
+ 4.292000000e-07 V_hig
+ 4.292010000e-07 V_hig
+ 4.293000000e-07 V_hig
+ 4.293010000e-07 V_hig
+ 4.294000000e-07 V_hig
+ 4.294010000e-07 V_hig
+ 4.295000000e-07 V_hig
+ 4.295010000e-07 V_hig
+ 4.296000000e-07 V_hig
+ 4.296010000e-07 V_hig
+ 4.297000000e-07 V_hig
+ 4.297010000e-07 V_hig
+ 4.298000000e-07 V_hig
+ 4.298010000e-07 V_hig
+ 4.299000000e-07 V_hig
+ 4.299010000e-07 V_hig
+ 4.300000000e-07 V_hig
+ 4.300010000e-07 V_hig
+ 4.301000000e-07 V_hig
+ 4.301010000e-07 V_hig
+ 4.302000000e-07 V_hig
+ 4.302010000e-07 V_hig
+ 4.303000000e-07 V_hig
+ 4.303010000e-07 V_hig
+ 4.304000000e-07 V_hig
+ 4.304010000e-07 V_hig
+ 4.305000000e-07 V_hig
+ 4.305010000e-07 V_hig
+ 4.306000000e-07 V_hig
+ 4.306010000e-07 V_hig
+ 4.307000000e-07 V_hig
+ 4.307010000e-07 V_hig
+ 4.308000000e-07 V_hig
+ 4.308010000e-07 V_hig
+ 4.309000000e-07 V_hig
+ 4.309010000e-07 V_hig
+ 4.310000000e-07 V_hig
+ 4.310010000e-07 V_hig
+ 4.311000000e-07 V_hig
+ 4.311010000e-07 V_hig
+ 4.312000000e-07 V_hig
+ 4.312010000e-07 V_hig
+ 4.313000000e-07 V_hig
+ 4.313010000e-07 V_hig
+ 4.314000000e-07 V_hig
+ 4.314010000e-07 V_hig
+ 4.315000000e-07 V_hig
+ 4.315010000e-07 V_hig
+ 4.316000000e-07 V_hig
+ 4.316010000e-07 V_hig
+ 4.317000000e-07 V_hig
+ 4.317010000e-07 V_hig
+ 4.318000000e-07 V_hig
+ 4.318010000e-07 V_hig
+ 4.319000000e-07 V_hig
+ 4.319010000e-07 V_low
+ 4.320000000e-07 V_low
+ 4.320010000e-07 V_low
+ 4.321000000e-07 V_low
+ 4.321010000e-07 V_low
+ 4.322000000e-07 V_low
+ 4.322010000e-07 V_low
+ 4.323000000e-07 V_low
+ 4.323010000e-07 V_low
+ 4.324000000e-07 V_low
+ 4.324010000e-07 V_low
+ 4.325000000e-07 V_low
+ 4.325010000e-07 V_low
+ 4.326000000e-07 V_low
+ 4.326010000e-07 V_low
+ 4.327000000e-07 V_low
+ 4.327010000e-07 V_low
+ 4.328000000e-07 V_low
+ 4.328010000e-07 V_low
+ 4.329000000e-07 V_low
+ 4.329010000e-07 V_low
+ 4.330000000e-07 V_low
+ 4.330010000e-07 V_low
+ 4.331000000e-07 V_low
+ 4.331010000e-07 V_low
+ 4.332000000e-07 V_low
+ 4.332010000e-07 V_low
+ 4.333000000e-07 V_low
+ 4.333010000e-07 V_low
+ 4.334000000e-07 V_low
+ 4.334010000e-07 V_low
+ 4.335000000e-07 V_low
+ 4.335010000e-07 V_low
+ 4.336000000e-07 V_low
+ 4.336010000e-07 V_low
+ 4.337000000e-07 V_low
+ 4.337010000e-07 V_low
+ 4.338000000e-07 V_low
+ 4.338010000e-07 V_low
+ 4.339000000e-07 V_low
+ 4.339010000e-07 V_hig
+ 4.340000000e-07 V_hig
+ 4.340010000e-07 V_hig
+ 4.341000000e-07 V_hig
+ 4.341010000e-07 V_hig
+ 4.342000000e-07 V_hig
+ 4.342010000e-07 V_hig
+ 4.343000000e-07 V_hig
+ 4.343010000e-07 V_hig
+ 4.344000000e-07 V_hig
+ 4.344010000e-07 V_hig
+ 4.345000000e-07 V_hig
+ 4.345010000e-07 V_hig
+ 4.346000000e-07 V_hig
+ 4.346010000e-07 V_hig
+ 4.347000000e-07 V_hig
+ 4.347010000e-07 V_hig
+ 4.348000000e-07 V_hig
+ 4.348010000e-07 V_hig
+ 4.349000000e-07 V_hig
+ 4.349010000e-07 V_hig
+ 4.350000000e-07 V_hig
+ 4.350010000e-07 V_hig
+ 4.351000000e-07 V_hig
+ 4.351010000e-07 V_hig
+ 4.352000000e-07 V_hig
+ 4.352010000e-07 V_hig
+ 4.353000000e-07 V_hig
+ 4.353010000e-07 V_hig
+ 4.354000000e-07 V_hig
+ 4.354010000e-07 V_hig
+ 4.355000000e-07 V_hig
+ 4.355010000e-07 V_hig
+ 4.356000000e-07 V_hig
+ 4.356010000e-07 V_hig
+ 4.357000000e-07 V_hig
+ 4.357010000e-07 V_hig
+ 4.358000000e-07 V_hig
+ 4.358010000e-07 V_hig
+ 4.359000000e-07 V_hig
+ 4.359010000e-07 V_hig
+ 4.360000000e-07 V_hig
+ 4.360010000e-07 V_hig
+ 4.361000000e-07 V_hig
+ 4.361010000e-07 V_hig
+ 4.362000000e-07 V_hig
+ 4.362010000e-07 V_hig
+ 4.363000000e-07 V_hig
+ 4.363010000e-07 V_hig
+ 4.364000000e-07 V_hig
+ 4.364010000e-07 V_hig
+ 4.365000000e-07 V_hig
+ 4.365010000e-07 V_hig
+ 4.366000000e-07 V_hig
+ 4.366010000e-07 V_hig
+ 4.367000000e-07 V_hig
+ 4.367010000e-07 V_hig
+ 4.368000000e-07 V_hig
+ 4.368010000e-07 V_hig
+ 4.369000000e-07 V_hig
+ 4.369010000e-07 V_hig
+ 4.370000000e-07 V_hig
+ 4.370010000e-07 V_hig
+ 4.371000000e-07 V_hig
+ 4.371010000e-07 V_hig
+ 4.372000000e-07 V_hig
+ 4.372010000e-07 V_hig
+ 4.373000000e-07 V_hig
+ 4.373010000e-07 V_hig
+ 4.374000000e-07 V_hig
+ 4.374010000e-07 V_hig
+ 4.375000000e-07 V_hig
+ 4.375010000e-07 V_hig
+ 4.376000000e-07 V_hig
+ 4.376010000e-07 V_hig
+ 4.377000000e-07 V_hig
+ 4.377010000e-07 V_hig
+ 4.378000000e-07 V_hig
+ 4.378010000e-07 V_hig
+ 4.379000000e-07 V_hig
+ 4.379010000e-07 V_hig
+ 4.380000000e-07 V_hig
+ 4.380010000e-07 V_hig
+ 4.381000000e-07 V_hig
+ 4.381010000e-07 V_hig
+ 4.382000000e-07 V_hig
+ 4.382010000e-07 V_hig
+ 4.383000000e-07 V_hig
+ 4.383010000e-07 V_hig
+ 4.384000000e-07 V_hig
+ 4.384010000e-07 V_hig
+ 4.385000000e-07 V_hig
+ 4.385010000e-07 V_hig
+ 4.386000000e-07 V_hig
+ 4.386010000e-07 V_hig
+ 4.387000000e-07 V_hig
+ 4.387010000e-07 V_hig
+ 4.388000000e-07 V_hig
+ 4.388010000e-07 V_hig
+ 4.389000000e-07 V_hig
+ 4.389010000e-07 V_hig
+ 4.390000000e-07 V_hig
+ 4.390010000e-07 V_hig
+ 4.391000000e-07 V_hig
+ 4.391010000e-07 V_hig
+ 4.392000000e-07 V_hig
+ 4.392010000e-07 V_hig
+ 4.393000000e-07 V_hig
+ 4.393010000e-07 V_hig
+ 4.394000000e-07 V_hig
+ 4.394010000e-07 V_hig
+ 4.395000000e-07 V_hig
+ 4.395010000e-07 V_hig
+ 4.396000000e-07 V_hig
+ 4.396010000e-07 V_hig
+ 4.397000000e-07 V_hig
+ 4.397010000e-07 V_hig
+ 4.398000000e-07 V_hig
+ 4.398010000e-07 V_hig
+ 4.399000000e-07 V_hig
+ 4.399010000e-07 V_low
+ 4.400000000e-07 V_low
+ 4.400010000e-07 V_low
+ 4.401000000e-07 V_low
+ 4.401010000e-07 V_low
+ 4.402000000e-07 V_low
+ 4.402010000e-07 V_low
+ 4.403000000e-07 V_low
+ 4.403010000e-07 V_low
+ 4.404000000e-07 V_low
+ 4.404010000e-07 V_low
+ 4.405000000e-07 V_low
+ 4.405010000e-07 V_low
+ 4.406000000e-07 V_low
+ 4.406010000e-07 V_low
+ 4.407000000e-07 V_low
+ 4.407010000e-07 V_low
+ 4.408000000e-07 V_low
+ 4.408010000e-07 V_low
+ 4.409000000e-07 V_low
+ 4.409010000e-07 V_low
+ 4.410000000e-07 V_low
+ 4.410010000e-07 V_low
+ 4.411000000e-07 V_low
+ 4.411010000e-07 V_low
+ 4.412000000e-07 V_low
+ 4.412010000e-07 V_low
+ 4.413000000e-07 V_low
+ 4.413010000e-07 V_low
+ 4.414000000e-07 V_low
+ 4.414010000e-07 V_low
+ 4.415000000e-07 V_low
+ 4.415010000e-07 V_low
+ 4.416000000e-07 V_low
+ 4.416010000e-07 V_low
+ 4.417000000e-07 V_low
+ 4.417010000e-07 V_low
+ 4.418000000e-07 V_low
+ 4.418010000e-07 V_low
+ 4.419000000e-07 V_low
+ 4.419010000e-07 V_hig
+ 4.420000000e-07 V_hig
+ 4.420010000e-07 V_hig
+ 4.421000000e-07 V_hig
+ 4.421010000e-07 V_hig
+ 4.422000000e-07 V_hig
+ 4.422010000e-07 V_hig
+ 4.423000000e-07 V_hig
+ 4.423010000e-07 V_hig
+ 4.424000000e-07 V_hig
+ 4.424010000e-07 V_hig
+ 4.425000000e-07 V_hig
+ 4.425010000e-07 V_hig
+ 4.426000000e-07 V_hig
+ 4.426010000e-07 V_hig
+ 4.427000000e-07 V_hig
+ 4.427010000e-07 V_hig
+ 4.428000000e-07 V_hig
+ 4.428010000e-07 V_hig
+ 4.429000000e-07 V_hig
+ 4.429010000e-07 V_low
+ 4.430000000e-07 V_low
+ 4.430010000e-07 V_low
+ 4.431000000e-07 V_low
+ 4.431010000e-07 V_low
+ 4.432000000e-07 V_low
+ 4.432010000e-07 V_low
+ 4.433000000e-07 V_low
+ 4.433010000e-07 V_low
+ 4.434000000e-07 V_low
+ 4.434010000e-07 V_low
+ 4.435000000e-07 V_low
+ 4.435010000e-07 V_low
+ 4.436000000e-07 V_low
+ 4.436010000e-07 V_low
+ 4.437000000e-07 V_low
+ 4.437010000e-07 V_low
+ 4.438000000e-07 V_low
+ 4.438010000e-07 V_low
+ 4.439000000e-07 V_low
+ 4.439010000e-07 V_low
+ 4.440000000e-07 V_low
+ 4.440010000e-07 V_low
+ 4.441000000e-07 V_low
+ 4.441010000e-07 V_low
+ 4.442000000e-07 V_low
+ 4.442010000e-07 V_low
+ 4.443000000e-07 V_low
+ 4.443010000e-07 V_low
+ 4.444000000e-07 V_low
+ 4.444010000e-07 V_low
+ 4.445000000e-07 V_low
+ 4.445010000e-07 V_low
+ 4.446000000e-07 V_low
+ 4.446010000e-07 V_low
+ 4.447000000e-07 V_low
+ 4.447010000e-07 V_low
+ 4.448000000e-07 V_low
+ 4.448010000e-07 V_low
+ 4.449000000e-07 V_low
+ 4.449010000e-07 V_low
+ 4.450000000e-07 V_low
+ 4.450010000e-07 V_low
+ 4.451000000e-07 V_low
+ 4.451010000e-07 V_low
+ 4.452000000e-07 V_low
+ 4.452010000e-07 V_low
+ 4.453000000e-07 V_low
+ 4.453010000e-07 V_low
+ 4.454000000e-07 V_low
+ 4.454010000e-07 V_low
+ 4.455000000e-07 V_low
+ 4.455010000e-07 V_low
+ 4.456000000e-07 V_low
+ 4.456010000e-07 V_low
+ 4.457000000e-07 V_low
+ 4.457010000e-07 V_low
+ 4.458000000e-07 V_low
+ 4.458010000e-07 V_low
+ 4.459000000e-07 V_low
+ 4.459010000e-07 V_low
+ 4.460000000e-07 V_low
+ 4.460010000e-07 V_low
+ 4.461000000e-07 V_low
+ 4.461010000e-07 V_low
+ 4.462000000e-07 V_low
+ 4.462010000e-07 V_low
+ 4.463000000e-07 V_low
+ 4.463010000e-07 V_low
+ 4.464000000e-07 V_low
+ 4.464010000e-07 V_low
+ 4.465000000e-07 V_low
+ 4.465010000e-07 V_low
+ 4.466000000e-07 V_low
+ 4.466010000e-07 V_low
+ 4.467000000e-07 V_low
+ 4.467010000e-07 V_low
+ 4.468000000e-07 V_low
+ 4.468010000e-07 V_low
+ 4.469000000e-07 V_low
+ 4.469010000e-07 V_hig
+ 4.470000000e-07 V_hig
+ 4.470010000e-07 V_hig
+ 4.471000000e-07 V_hig
+ 4.471010000e-07 V_hig
+ 4.472000000e-07 V_hig
+ 4.472010000e-07 V_hig
+ 4.473000000e-07 V_hig
+ 4.473010000e-07 V_hig
+ 4.474000000e-07 V_hig
+ 4.474010000e-07 V_hig
+ 4.475000000e-07 V_hig
+ 4.475010000e-07 V_hig
+ 4.476000000e-07 V_hig
+ 4.476010000e-07 V_hig
+ 4.477000000e-07 V_hig
+ 4.477010000e-07 V_hig
+ 4.478000000e-07 V_hig
+ 4.478010000e-07 V_hig
+ 4.479000000e-07 V_hig
+ 4.479010000e-07 V_low
+ 4.480000000e-07 V_low
+ 4.480010000e-07 V_low
+ 4.481000000e-07 V_low
+ 4.481010000e-07 V_low
+ 4.482000000e-07 V_low
+ 4.482010000e-07 V_low
+ 4.483000000e-07 V_low
+ 4.483010000e-07 V_low
+ 4.484000000e-07 V_low
+ 4.484010000e-07 V_low
+ 4.485000000e-07 V_low
+ 4.485010000e-07 V_low
+ 4.486000000e-07 V_low
+ 4.486010000e-07 V_low
+ 4.487000000e-07 V_low
+ 4.487010000e-07 V_low
+ 4.488000000e-07 V_low
+ 4.488010000e-07 V_low
+ 4.489000000e-07 V_low
+ 4.489010000e-07 V_hig
+ 4.490000000e-07 V_hig
+ 4.490010000e-07 V_hig
+ 4.491000000e-07 V_hig
+ 4.491010000e-07 V_hig
+ 4.492000000e-07 V_hig
+ 4.492010000e-07 V_hig
+ 4.493000000e-07 V_hig
+ 4.493010000e-07 V_hig
+ 4.494000000e-07 V_hig
+ 4.494010000e-07 V_hig
+ 4.495000000e-07 V_hig
+ 4.495010000e-07 V_hig
+ 4.496000000e-07 V_hig
+ 4.496010000e-07 V_hig
+ 4.497000000e-07 V_hig
+ 4.497010000e-07 V_hig
+ 4.498000000e-07 V_hig
+ 4.498010000e-07 V_hig
+ 4.499000000e-07 V_hig
+ 4.499010000e-07 V_hig
+ 4.500000000e-07 V_hig
+ 4.500010000e-07 V_hig
+ 4.501000000e-07 V_hig
+ 4.501010000e-07 V_hig
+ 4.502000000e-07 V_hig
+ 4.502010000e-07 V_hig
+ 4.503000000e-07 V_hig
+ 4.503010000e-07 V_hig
+ 4.504000000e-07 V_hig
+ 4.504010000e-07 V_hig
+ 4.505000000e-07 V_hig
+ 4.505010000e-07 V_hig
+ 4.506000000e-07 V_hig
+ 4.506010000e-07 V_hig
+ 4.507000000e-07 V_hig
+ 4.507010000e-07 V_hig
+ 4.508000000e-07 V_hig
+ 4.508010000e-07 V_hig
+ 4.509000000e-07 V_hig
+ 4.509010000e-07 V_hig
+ 4.510000000e-07 V_hig
+ 4.510010000e-07 V_hig
+ 4.511000000e-07 V_hig
+ 4.511010000e-07 V_hig
+ 4.512000000e-07 V_hig
+ 4.512010000e-07 V_hig
+ 4.513000000e-07 V_hig
+ 4.513010000e-07 V_hig
+ 4.514000000e-07 V_hig
+ 4.514010000e-07 V_hig
+ 4.515000000e-07 V_hig
+ 4.515010000e-07 V_hig
+ 4.516000000e-07 V_hig
+ 4.516010000e-07 V_hig
+ 4.517000000e-07 V_hig
+ 4.517010000e-07 V_hig
+ 4.518000000e-07 V_hig
+ 4.518010000e-07 V_hig
+ 4.519000000e-07 V_hig
+ 4.519010000e-07 V_hig
+ 4.520000000e-07 V_hig
+ 4.520010000e-07 V_hig
+ 4.521000000e-07 V_hig
+ 4.521010000e-07 V_hig
+ 4.522000000e-07 V_hig
+ 4.522010000e-07 V_hig
+ 4.523000000e-07 V_hig
+ 4.523010000e-07 V_hig
+ 4.524000000e-07 V_hig
+ 4.524010000e-07 V_hig
+ 4.525000000e-07 V_hig
+ 4.525010000e-07 V_hig
+ 4.526000000e-07 V_hig
+ 4.526010000e-07 V_hig
+ 4.527000000e-07 V_hig
+ 4.527010000e-07 V_hig
+ 4.528000000e-07 V_hig
+ 4.528010000e-07 V_hig
+ 4.529000000e-07 V_hig
+ 4.529010000e-07 V_low
+ 4.530000000e-07 V_low
+ 4.530010000e-07 V_low
+ 4.531000000e-07 V_low
+ 4.531010000e-07 V_low
+ 4.532000000e-07 V_low
+ 4.532010000e-07 V_low
+ 4.533000000e-07 V_low
+ 4.533010000e-07 V_low
+ 4.534000000e-07 V_low
+ 4.534010000e-07 V_low
+ 4.535000000e-07 V_low
+ 4.535010000e-07 V_low
+ 4.536000000e-07 V_low
+ 4.536010000e-07 V_low
+ 4.537000000e-07 V_low
+ 4.537010000e-07 V_low
+ 4.538000000e-07 V_low
+ 4.538010000e-07 V_low
+ 4.539000000e-07 V_low
+ 4.539010000e-07 V_low
+ 4.540000000e-07 V_low
+ 4.540010000e-07 V_low
+ 4.541000000e-07 V_low
+ 4.541010000e-07 V_low
+ 4.542000000e-07 V_low
+ 4.542010000e-07 V_low
+ 4.543000000e-07 V_low
+ 4.543010000e-07 V_low
+ 4.544000000e-07 V_low
+ 4.544010000e-07 V_low
+ 4.545000000e-07 V_low
+ 4.545010000e-07 V_low
+ 4.546000000e-07 V_low
+ 4.546010000e-07 V_low
+ 4.547000000e-07 V_low
+ 4.547010000e-07 V_low
+ 4.548000000e-07 V_low
+ 4.548010000e-07 V_low
+ 4.549000000e-07 V_low
+ 4.549010000e-07 V_low
+ 4.550000000e-07 V_low
+ 4.550010000e-07 V_low
+ 4.551000000e-07 V_low
+ 4.551010000e-07 V_low
+ 4.552000000e-07 V_low
+ 4.552010000e-07 V_low
+ 4.553000000e-07 V_low
+ 4.553010000e-07 V_low
+ 4.554000000e-07 V_low
+ 4.554010000e-07 V_low
+ 4.555000000e-07 V_low
+ 4.555010000e-07 V_low
+ 4.556000000e-07 V_low
+ 4.556010000e-07 V_low
+ 4.557000000e-07 V_low
+ 4.557010000e-07 V_low
+ 4.558000000e-07 V_low
+ 4.558010000e-07 V_low
+ 4.559000000e-07 V_low
+ 4.559010000e-07 V_low
+ 4.560000000e-07 V_low
+ 4.560010000e-07 V_low
+ 4.561000000e-07 V_low
+ 4.561010000e-07 V_low
+ 4.562000000e-07 V_low
+ 4.562010000e-07 V_low
+ 4.563000000e-07 V_low
+ 4.563010000e-07 V_low
+ 4.564000000e-07 V_low
+ 4.564010000e-07 V_low
+ 4.565000000e-07 V_low
+ 4.565010000e-07 V_low
+ 4.566000000e-07 V_low
+ 4.566010000e-07 V_low
+ 4.567000000e-07 V_low
+ 4.567010000e-07 V_low
+ 4.568000000e-07 V_low
+ 4.568010000e-07 V_low
+ 4.569000000e-07 V_low
+ 4.569010000e-07 V_low
+ 4.570000000e-07 V_low
+ 4.570010000e-07 V_low
+ 4.571000000e-07 V_low
+ 4.571010000e-07 V_low
+ 4.572000000e-07 V_low
+ 4.572010000e-07 V_low
+ 4.573000000e-07 V_low
+ 4.573010000e-07 V_low
+ 4.574000000e-07 V_low
+ 4.574010000e-07 V_low
+ 4.575000000e-07 V_low
+ 4.575010000e-07 V_low
+ 4.576000000e-07 V_low
+ 4.576010000e-07 V_low
+ 4.577000000e-07 V_low
+ 4.577010000e-07 V_low
+ 4.578000000e-07 V_low
+ 4.578010000e-07 V_low
+ 4.579000000e-07 V_low
+ 4.579010000e-07 V_low
+ 4.580000000e-07 V_low
+ 4.580010000e-07 V_low
+ 4.581000000e-07 V_low
+ 4.581010000e-07 V_low
+ 4.582000000e-07 V_low
+ 4.582010000e-07 V_low
+ 4.583000000e-07 V_low
+ 4.583010000e-07 V_low
+ 4.584000000e-07 V_low
+ 4.584010000e-07 V_low
+ 4.585000000e-07 V_low
+ 4.585010000e-07 V_low
+ 4.586000000e-07 V_low
+ 4.586010000e-07 V_low
+ 4.587000000e-07 V_low
+ 4.587010000e-07 V_low
+ 4.588000000e-07 V_low
+ 4.588010000e-07 V_low
+ 4.589000000e-07 V_low
+ 4.589010000e-07 V_low
+ 4.590000000e-07 V_low
+ 4.590010000e-07 V_low
+ 4.591000000e-07 V_low
+ 4.591010000e-07 V_low
+ 4.592000000e-07 V_low
+ 4.592010000e-07 V_low
+ 4.593000000e-07 V_low
+ 4.593010000e-07 V_low
+ 4.594000000e-07 V_low
+ 4.594010000e-07 V_low
+ 4.595000000e-07 V_low
+ 4.595010000e-07 V_low
+ 4.596000000e-07 V_low
+ 4.596010000e-07 V_low
+ 4.597000000e-07 V_low
+ 4.597010000e-07 V_low
+ 4.598000000e-07 V_low
+ 4.598010000e-07 V_low
+ 4.599000000e-07 V_low
+ 4.599010000e-07 V_low
+ 4.600000000e-07 V_low
+ 4.600010000e-07 V_low
+ 4.601000000e-07 V_low
+ 4.601010000e-07 V_low
+ 4.602000000e-07 V_low
+ 4.602010000e-07 V_low
+ 4.603000000e-07 V_low
+ 4.603010000e-07 V_low
+ 4.604000000e-07 V_low
+ 4.604010000e-07 V_low
+ 4.605000000e-07 V_low
+ 4.605010000e-07 V_low
+ 4.606000000e-07 V_low
+ 4.606010000e-07 V_low
+ 4.607000000e-07 V_low
+ 4.607010000e-07 V_low
+ 4.608000000e-07 V_low
+ 4.608010000e-07 V_low
+ 4.609000000e-07 V_low
+ 4.609010000e-07 V_low
+ 4.610000000e-07 V_low
+ 4.610010000e-07 V_low
+ 4.611000000e-07 V_low
+ 4.611010000e-07 V_low
+ 4.612000000e-07 V_low
+ 4.612010000e-07 V_low
+ 4.613000000e-07 V_low
+ 4.613010000e-07 V_low
+ 4.614000000e-07 V_low
+ 4.614010000e-07 V_low
+ 4.615000000e-07 V_low
+ 4.615010000e-07 V_low
+ 4.616000000e-07 V_low
+ 4.616010000e-07 V_low
+ 4.617000000e-07 V_low
+ 4.617010000e-07 V_low
+ 4.618000000e-07 V_low
+ 4.618010000e-07 V_low
+ 4.619000000e-07 V_low
+ 4.619010000e-07 V_hig
+ 4.620000000e-07 V_hig
+ 4.620010000e-07 V_hig
+ 4.621000000e-07 V_hig
+ 4.621010000e-07 V_hig
+ 4.622000000e-07 V_hig
+ 4.622010000e-07 V_hig
+ 4.623000000e-07 V_hig
+ 4.623010000e-07 V_hig
+ 4.624000000e-07 V_hig
+ 4.624010000e-07 V_hig
+ 4.625000000e-07 V_hig
+ 4.625010000e-07 V_hig
+ 4.626000000e-07 V_hig
+ 4.626010000e-07 V_hig
+ 4.627000000e-07 V_hig
+ 4.627010000e-07 V_hig
+ 4.628000000e-07 V_hig
+ 4.628010000e-07 V_hig
+ 4.629000000e-07 V_hig
+ 4.629010000e-07 V_hig
+ 4.630000000e-07 V_hig
+ 4.630010000e-07 V_hig
+ 4.631000000e-07 V_hig
+ 4.631010000e-07 V_hig
+ 4.632000000e-07 V_hig
+ 4.632010000e-07 V_hig
+ 4.633000000e-07 V_hig
+ 4.633010000e-07 V_hig
+ 4.634000000e-07 V_hig
+ 4.634010000e-07 V_hig
+ 4.635000000e-07 V_hig
+ 4.635010000e-07 V_hig
+ 4.636000000e-07 V_hig
+ 4.636010000e-07 V_hig
+ 4.637000000e-07 V_hig
+ 4.637010000e-07 V_hig
+ 4.638000000e-07 V_hig
+ 4.638010000e-07 V_hig
+ 4.639000000e-07 V_hig
+ 4.639010000e-07 V_hig
+ 4.640000000e-07 V_hig
+ 4.640010000e-07 V_hig
+ 4.641000000e-07 V_hig
+ 4.641010000e-07 V_hig
+ 4.642000000e-07 V_hig
+ 4.642010000e-07 V_hig
+ 4.643000000e-07 V_hig
+ 4.643010000e-07 V_hig
+ 4.644000000e-07 V_hig
+ 4.644010000e-07 V_hig
+ 4.645000000e-07 V_hig
+ 4.645010000e-07 V_hig
+ 4.646000000e-07 V_hig
+ 4.646010000e-07 V_hig
+ 4.647000000e-07 V_hig
+ 4.647010000e-07 V_hig
+ 4.648000000e-07 V_hig
+ 4.648010000e-07 V_hig
+ 4.649000000e-07 V_hig
+ 4.649010000e-07 V_low
+ 4.650000000e-07 V_low
+ 4.650010000e-07 V_low
+ 4.651000000e-07 V_low
+ 4.651010000e-07 V_low
+ 4.652000000e-07 V_low
+ 4.652010000e-07 V_low
+ 4.653000000e-07 V_low
+ 4.653010000e-07 V_low
+ 4.654000000e-07 V_low
+ 4.654010000e-07 V_low
+ 4.655000000e-07 V_low
+ 4.655010000e-07 V_low
+ 4.656000000e-07 V_low
+ 4.656010000e-07 V_low
+ 4.657000000e-07 V_low
+ 4.657010000e-07 V_low
+ 4.658000000e-07 V_low
+ 4.658010000e-07 V_low
+ 4.659000000e-07 V_low
+ 4.659010000e-07 V_low
+ 4.660000000e-07 V_low
+ 4.660010000e-07 V_low
+ 4.661000000e-07 V_low
+ 4.661010000e-07 V_low
+ 4.662000000e-07 V_low
+ 4.662010000e-07 V_low
+ 4.663000000e-07 V_low
+ 4.663010000e-07 V_low
+ 4.664000000e-07 V_low
+ 4.664010000e-07 V_low
+ 4.665000000e-07 V_low
+ 4.665010000e-07 V_low
+ 4.666000000e-07 V_low
+ 4.666010000e-07 V_low
+ 4.667000000e-07 V_low
+ 4.667010000e-07 V_low
+ 4.668000000e-07 V_low
+ 4.668010000e-07 V_low
+ 4.669000000e-07 V_low
+ 4.669010000e-07 V_low
+ 4.670000000e-07 V_low
+ 4.670010000e-07 V_low
+ 4.671000000e-07 V_low
+ 4.671010000e-07 V_low
+ 4.672000000e-07 V_low
+ 4.672010000e-07 V_low
+ 4.673000000e-07 V_low
+ 4.673010000e-07 V_low
+ 4.674000000e-07 V_low
+ 4.674010000e-07 V_low
+ 4.675000000e-07 V_low
+ 4.675010000e-07 V_low
+ 4.676000000e-07 V_low
+ 4.676010000e-07 V_low
+ 4.677000000e-07 V_low
+ 4.677010000e-07 V_low
+ 4.678000000e-07 V_low
+ 4.678010000e-07 V_low
+ 4.679000000e-07 V_low
+ 4.679010000e-07 V_low
+ 4.680000000e-07 V_low
+ 4.680010000e-07 V_low
+ 4.681000000e-07 V_low
+ 4.681010000e-07 V_low
+ 4.682000000e-07 V_low
+ 4.682010000e-07 V_low
+ 4.683000000e-07 V_low
+ 4.683010000e-07 V_low
+ 4.684000000e-07 V_low
+ 4.684010000e-07 V_low
+ 4.685000000e-07 V_low
+ 4.685010000e-07 V_low
+ 4.686000000e-07 V_low
+ 4.686010000e-07 V_low
+ 4.687000000e-07 V_low
+ 4.687010000e-07 V_low
+ 4.688000000e-07 V_low
+ 4.688010000e-07 V_low
+ 4.689000000e-07 V_low
+ 4.689010000e-07 V_hig
+ 4.690000000e-07 V_hig
+ 4.690010000e-07 V_hig
+ 4.691000000e-07 V_hig
+ 4.691010000e-07 V_hig
+ 4.692000000e-07 V_hig
+ 4.692010000e-07 V_hig
+ 4.693000000e-07 V_hig
+ 4.693010000e-07 V_hig
+ 4.694000000e-07 V_hig
+ 4.694010000e-07 V_hig
+ 4.695000000e-07 V_hig
+ 4.695010000e-07 V_hig
+ 4.696000000e-07 V_hig
+ 4.696010000e-07 V_hig
+ 4.697000000e-07 V_hig
+ 4.697010000e-07 V_hig
+ 4.698000000e-07 V_hig
+ 4.698010000e-07 V_hig
+ 4.699000000e-07 V_hig
+ 4.699010000e-07 V_low
+ 4.700000000e-07 V_low
+ 4.700010000e-07 V_low
+ 4.701000000e-07 V_low
+ 4.701010000e-07 V_low
+ 4.702000000e-07 V_low
+ 4.702010000e-07 V_low
+ 4.703000000e-07 V_low
+ 4.703010000e-07 V_low
+ 4.704000000e-07 V_low
+ 4.704010000e-07 V_low
+ 4.705000000e-07 V_low
+ 4.705010000e-07 V_low
+ 4.706000000e-07 V_low
+ 4.706010000e-07 V_low
+ 4.707000000e-07 V_low
+ 4.707010000e-07 V_low
+ 4.708000000e-07 V_low
+ 4.708010000e-07 V_low
+ 4.709000000e-07 V_low
+ 4.709010000e-07 V_low
+ 4.710000000e-07 V_low
+ 4.710010000e-07 V_low
+ 4.711000000e-07 V_low
+ 4.711010000e-07 V_low
+ 4.712000000e-07 V_low
+ 4.712010000e-07 V_low
+ 4.713000000e-07 V_low
+ 4.713010000e-07 V_low
+ 4.714000000e-07 V_low
+ 4.714010000e-07 V_low
+ 4.715000000e-07 V_low
+ 4.715010000e-07 V_low
+ 4.716000000e-07 V_low
+ 4.716010000e-07 V_low
+ 4.717000000e-07 V_low
+ 4.717010000e-07 V_low
+ 4.718000000e-07 V_low
+ 4.718010000e-07 V_low
+ 4.719000000e-07 V_low
+ 4.719010000e-07 V_low
+ 4.720000000e-07 V_low
+ 4.720010000e-07 V_low
+ 4.721000000e-07 V_low
+ 4.721010000e-07 V_low
+ 4.722000000e-07 V_low
+ 4.722010000e-07 V_low
+ 4.723000000e-07 V_low
+ 4.723010000e-07 V_low
+ 4.724000000e-07 V_low
+ 4.724010000e-07 V_low
+ 4.725000000e-07 V_low
+ 4.725010000e-07 V_low
+ 4.726000000e-07 V_low
+ 4.726010000e-07 V_low
+ 4.727000000e-07 V_low
+ 4.727010000e-07 V_low
+ 4.728000000e-07 V_low
+ 4.728010000e-07 V_low
+ 4.729000000e-07 V_low
+ 4.729010000e-07 V_hig
+ 4.730000000e-07 V_hig
+ 4.730010000e-07 V_hig
+ 4.731000000e-07 V_hig
+ 4.731010000e-07 V_hig
+ 4.732000000e-07 V_hig
+ 4.732010000e-07 V_hig
+ 4.733000000e-07 V_hig
+ 4.733010000e-07 V_hig
+ 4.734000000e-07 V_hig
+ 4.734010000e-07 V_hig
+ 4.735000000e-07 V_hig
+ 4.735010000e-07 V_hig
+ 4.736000000e-07 V_hig
+ 4.736010000e-07 V_hig
+ 4.737000000e-07 V_hig
+ 4.737010000e-07 V_hig
+ 4.738000000e-07 V_hig
+ 4.738010000e-07 V_hig
+ 4.739000000e-07 V_hig
+ 4.739010000e-07 V_low
+ 4.740000000e-07 V_low
+ 4.740010000e-07 V_low
+ 4.741000000e-07 V_low
+ 4.741010000e-07 V_low
+ 4.742000000e-07 V_low
+ 4.742010000e-07 V_low
+ 4.743000000e-07 V_low
+ 4.743010000e-07 V_low
+ 4.744000000e-07 V_low
+ 4.744010000e-07 V_low
+ 4.745000000e-07 V_low
+ 4.745010000e-07 V_low
+ 4.746000000e-07 V_low
+ 4.746010000e-07 V_low
+ 4.747000000e-07 V_low
+ 4.747010000e-07 V_low
+ 4.748000000e-07 V_low
+ 4.748010000e-07 V_low
+ 4.749000000e-07 V_low
+ 4.749010000e-07 V_hig
+ 4.750000000e-07 V_hig
+ 4.750010000e-07 V_hig
+ 4.751000000e-07 V_hig
+ 4.751010000e-07 V_hig
+ 4.752000000e-07 V_hig
+ 4.752010000e-07 V_hig
+ 4.753000000e-07 V_hig
+ 4.753010000e-07 V_hig
+ 4.754000000e-07 V_hig
+ 4.754010000e-07 V_hig
+ 4.755000000e-07 V_hig
+ 4.755010000e-07 V_hig
+ 4.756000000e-07 V_hig
+ 4.756010000e-07 V_hig
+ 4.757000000e-07 V_hig
+ 4.757010000e-07 V_hig
+ 4.758000000e-07 V_hig
+ 4.758010000e-07 V_hig
+ 4.759000000e-07 V_hig
+ 4.759010000e-07 V_low
+ 4.760000000e-07 V_low
+ 4.760010000e-07 V_low
+ 4.761000000e-07 V_low
+ 4.761010000e-07 V_low
+ 4.762000000e-07 V_low
+ 4.762010000e-07 V_low
+ 4.763000000e-07 V_low
+ 4.763010000e-07 V_low
+ 4.764000000e-07 V_low
+ 4.764010000e-07 V_low
+ 4.765000000e-07 V_low
+ 4.765010000e-07 V_low
+ 4.766000000e-07 V_low
+ 4.766010000e-07 V_low
+ 4.767000000e-07 V_low
+ 4.767010000e-07 V_low
+ 4.768000000e-07 V_low
+ 4.768010000e-07 V_low
+ 4.769000000e-07 V_low
+ 4.769010000e-07 V_hig
+ 4.770000000e-07 V_hig
+ 4.770010000e-07 V_hig
+ 4.771000000e-07 V_hig
+ 4.771010000e-07 V_hig
+ 4.772000000e-07 V_hig
+ 4.772010000e-07 V_hig
+ 4.773000000e-07 V_hig
+ 4.773010000e-07 V_hig
+ 4.774000000e-07 V_hig
+ 4.774010000e-07 V_hig
+ 4.775000000e-07 V_hig
+ 4.775010000e-07 V_hig
+ 4.776000000e-07 V_hig
+ 4.776010000e-07 V_hig
+ 4.777000000e-07 V_hig
+ 4.777010000e-07 V_hig
+ 4.778000000e-07 V_hig
+ 4.778010000e-07 V_hig
+ 4.779000000e-07 V_hig
+ 4.779010000e-07 V_hig
+ 4.780000000e-07 V_hig
+ 4.780010000e-07 V_hig
+ 4.781000000e-07 V_hig
+ 4.781010000e-07 V_hig
+ 4.782000000e-07 V_hig
+ 4.782010000e-07 V_hig
+ 4.783000000e-07 V_hig
+ 4.783010000e-07 V_hig
+ 4.784000000e-07 V_hig
+ 4.784010000e-07 V_hig
+ 4.785000000e-07 V_hig
+ 4.785010000e-07 V_hig
+ 4.786000000e-07 V_hig
+ 4.786010000e-07 V_hig
+ 4.787000000e-07 V_hig
+ 4.787010000e-07 V_hig
+ 4.788000000e-07 V_hig
+ 4.788010000e-07 V_hig
+ 4.789000000e-07 V_hig
+ 4.789010000e-07 V_hig
+ 4.790000000e-07 V_hig
+ 4.790010000e-07 V_hig
+ 4.791000000e-07 V_hig
+ 4.791010000e-07 V_hig
+ 4.792000000e-07 V_hig
+ 4.792010000e-07 V_hig
+ 4.793000000e-07 V_hig
+ 4.793010000e-07 V_hig
+ 4.794000000e-07 V_hig
+ 4.794010000e-07 V_hig
+ 4.795000000e-07 V_hig
+ 4.795010000e-07 V_hig
+ 4.796000000e-07 V_hig
+ 4.796010000e-07 V_hig
+ 4.797000000e-07 V_hig
+ 4.797010000e-07 V_hig
+ 4.798000000e-07 V_hig
+ 4.798010000e-07 V_hig
+ 4.799000000e-07 V_hig
+ 4.799010000e-07 V_low
+ 4.800000000e-07 V_low
+ 4.800010000e-07 V_low
+ 4.801000000e-07 V_low
+ 4.801010000e-07 V_low
+ 4.802000000e-07 V_low
+ 4.802010000e-07 V_low
+ 4.803000000e-07 V_low
+ 4.803010000e-07 V_low
+ 4.804000000e-07 V_low
+ 4.804010000e-07 V_low
+ 4.805000000e-07 V_low
+ 4.805010000e-07 V_low
+ 4.806000000e-07 V_low
+ 4.806010000e-07 V_low
+ 4.807000000e-07 V_low
+ 4.807010000e-07 V_low
+ 4.808000000e-07 V_low
+ 4.808010000e-07 V_low
+ 4.809000000e-07 V_low
+ 4.809010000e-07 V_low
+ 4.810000000e-07 V_low
+ 4.810010000e-07 V_low
+ 4.811000000e-07 V_low
+ 4.811010000e-07 V_low
+ 4.812000000e-07 V_low
+ 4.812010000e-07 V_low
+ 4.813000000e-07 V_low
+ 4.813010000e-07 V_low
+ 4.814000000e-07 V_low
+ 4.814010000e-07 V_low
+ 4.815000000e-07 V_low
+ 4.815010000e-07 V_low
+ 4.816000000e-07 V_low
+ 4.816010000e-07 V_low
+ 4.817000000e-07 V_low
+ 4.817010000e-07 V_low
+ 4.818000000e-07 V_low
+ 4.818010000e-07 V_low
+ 4.819000000e-07 V_low
+ 4.819010000e-07 V_low
+ 4.820000000e-07 V_low
+ 4.820010000e-07 V_low
+ 4.821000000e-07 V_low
+ 4.821010000e-07 V_low
+ 4.822000000e-07 V_low
+ 4.822010000e-07 V_low
+ 4.823000000e-07 V_low
+ 4.823010000e-07 V_low
+ 4.824000000e-07 V_low
+ 4.824010000e-07 V_low
+ 4.825000000e-07 V_low
+ 4.825010000e-07 V_low
+ 4.826000000e-07 V_low
+ 4.826010000e-07 V_low
+ 4.827000000e-07 V_low
+ 4.827010000e-07 V_low
+ 4.828000000e-07 V_low
+ 4.828010000e-07 V_low
+ 4.829000000e-07 V_low
+ 4.829010000e-07 V_low
+ 4.830000000e-07 V_low
+ 4.830010000e-07 V_low
+ 4.831000000e-07 V_low
+ 4.831010000e-07 V_low
+ 4.832000000e-07 V_low
+ 4.832010000e-07 V_low
+ 4.833000000e-07 V_low
+ 4.833010000e-07 V_low
+ 4.834000000e-07 V_low
+ 4.834010000e-07 V_low
+ 4.835000000e-07 V_low
+ 4.835010000e-07 V_low
+ 4.836000000e-07 V_low
+ 4.836010000e-07 V_low
+ 4.837000000e-07 V_low
+ 4.837010000e-07 V_low
+ 4.838000000e-07 V_low
+ 4.838010000e-07 V_low
+ 4.839000000e-07 V_low
+ 4.839010000e-07 V_low
+ 4.840000000e-07 V_low
+ 4.840010000e-07 V_low
+ 4.841000000e-07 V_low
+ 4.841010000e-07 V_low
+ 4.842000000e-07 V_low
+ 4.842010000e-07 V_low
+ 4.843000000e-07 V_low
+ 4.843010000e-07 V_low
+ 4.844000000e-07 V_low
+ 4.844010000e-07 V_low
+ 4.845000000e-07 V_low
+ 4.845010000e-07 V_low
+ 4.846000000e-07 V_low
+ 4.846010000e-07 V_low
+ 4.847000000e-07 V_low
+ 4.847010000e-07 V_low
+ 4.848000000e-07 V_low
+ 4.848010000e-07 V_low
+ 4.849000000e-07 V_low
+ 4.849010000e-07 V_low
+ 4.850000000e-07 V_low
+ 4.850010000e-07 V_low
+ 4.851000000e-07 V_low
+ 4.851010000e-07 V_low
+ 4.852000000e-07 V_low
+ 4.852010000e-07 V_low
+ 4.853000000e-07 V_low
+ 4.853010000e-07 V_low
+ 4.854000000e-07 V_low
+ 4.854010000e-07 V_low
+ 4.855000000e-07 V_low
+ 4.855010000e-07 V_low
+ 4.856000000e-07 V_low
+ 4.856010000e-07 V_low
+ 4.857000000e-07 V_low
+ 4.857010000e-07 V_low
+ 4.858000000e-07 V_low
+ 4.858010000e-07 V_low
+ 4.859000000e-07 V_low
+ 4.859010000e-07 V_hig
+ 4.860000000e-07 V_hig
+ 4.860010000e-07 V_hig
+ 4.861000000e-07 V_hig
+ 4.861010000e-07 V_hig
+ 4.862000000e-07 V_hig
+ 4.862010000e-07 V_hig
+ 4.863000000e-07 V_hig
+ 4.863010000e-07 V_hig
+ 4.864000000e-07 V_hig
+ 4.864010000e-07 V_hig
+ 4.865000000e-07 V_hig
+ 4.865010000e-07 V_hig
+ 4.866000000e-07 V_hig
+ 4.866010000e-07 V_hig
+ 4.867000000e-07 V_hig
+ 4.867010000e-07 V_hig
+ 4.868000000e-07 V_hig
+ 4.868010000e-07 V_hig
+ 4.869000000e-07 V_hig
+ 4.869010000e-07 V_low
+ 4.870000000e-07 V_low
+ 4.870010000e-07 V_low
+ 4.871000000e-07 V_low
+ 4.871010000e-07 V_low
+ 4.872000000e-07 V_low
+ 4.872010000e-07 V_low
+ 4.873000000e-07 V_low
+ 4.873010000e-07 V_low
+ 4.874000000e-07 V_low
+ 4.874010000e-07 V_low
+ 4.875000000e-07 V_low
+ 4.875010000e-07 V_low
+ 4.876000000e-07 V_low
+ 4.876010000e-07 V_low
+ 4.877000000e-07 V_low
+ 4.877010000e-07 V_low
+ 4.878000000e-07 V_low
+ 4.878010000e-07 V_low
+ 4.879000000e-07 V_low
+ 4.879010000e-07 V_low
+ 4.880000000e-07 V_low
+ 4.880010000e-07 V_low
+ 4.881000000e-07 V_low
+ 4.881010000e-07 V_low
+ 4.882000000e-07 V_low
+ 4.882010000e-07 V_low
+ 4.883000000e-07 V_low
+ 4.883010000e-07 V_low
+ 4.884000000e-07 V_low
+ 4.884010000e-07 V_low
+ 4.885000000e-07 V_low
+ 4.885010000e-07 V_low
+ 4.886000000e-07 V_low
+ 4.886010000e-07 V_low
+ 4.887000000e-07 V_low
+ 4.887010000e-07 V_low
+ 4.888000000e-07 V_low
+ 4.888010000e-07 V_low
+ 4.889000000e-07 V_low
+ 4.889010000e-07 V_hig
+ 4.890000000e-07 V_hig
+ 4.890010000e-07 V_hig
+ 4.891000000e-07 V_hig
+ 4.891010000e-07 V_hig
+ 4.892000000e-07 V_hig
+ 4.892010000e-07 V_hig
+ 4.893000000e-07 V_hig
+ 4.893010000e-07 V_hig
+ 4.894000000e-07 V_hig
+ 4.894010000e-07 V_hig
+ 4.895000000e-07 V_hig
+ 4.895010000e-07 V_hig
+ 4.896000000e-07 V_hig
+ 4.896010000e-07 V_hig
+ 4.897000000e-07 V_hig
+ 4.897010000e-07 V_hig
+ 4.898000000e-07 V_hig
+ 4.898010000e-07 V_hig
+ 4.899000000e-07 V_hig
+ 4.899010000e-07 V_hig
+ 4.900000000e-07 V_hig
+ 4.900010000e-07 V_hig
+ 4.901000000e-07 V_hig
+ 4.901010000e-07 V_hig
+ 4.902000000e-07 V_hig
+ 4.902010000e-07 V_hig
+ 4.903000000e-07 V_hig
+ 4.903010000e-07 V_hig
+ 4.904000000e-07 V_hig
+ 4.904010000e-07 V_hig
+ 4.905000000e-07 V_hig
+ 4.905010000e-07 V_hig
+ 4.906000000e-07 V_hig
+ 4.906010000e-07 V_hig
+ 4.907000000e-07 V_hig
+ 4.907010000e-07 V_hig
+ 4.908000000e-07 V_hig
+ 4.908010000e-07 V_hig
+ 4.909000000e-07 V_hig
+ 4.909010000e-07 V_hig
+ 4.910000000e-07 V_hig
+ 4.910010000e-07 V_hig
+ 4.911000000e-07 V_hig
+ 4.911010000e-07 V_hig
+ 4.912000000e-07 V_hig
+ 4.912010000e-07 V_hig
+ 4.913000000e-07 V_hig
+ 4.913010000e-07 V_hig
+ 4.914000000e-07 V_hig
+ 4.914010000e-07 V_hig
+ 4.915000000e-07 V_hig
+ 4.915010000e-07 V_hig
+ 4.916000000e-07 V_hig
+ 4.916010000e-07 V_hig
+ 4.917000000e-07 V_hig
+ 4.917010000e-07 V_hig
+ 4.918000000e-07 V_hig
+ 4.918010000e-07 V_hig
+ 4.919000000e-07 V_hig
+ 4.919010000e-07 V_low
+ 4.920000000e-07 V_low
+ 4.920010000e-07 V_low
+ 4.921000000e-07 V_low
+ 4.921010000e-07 V_low
+ 4.922000000e-07 V_low
+ 4.922010000e-07 V_low
+ 4.923000000e-07 V_low
+ 4.923010000e-07 V_low
+ 4.924000000e-07 V_low
+ 4.924010000e-07 V_low
+ 4.925000000e-07 V_low
+ 4.925010000e-07 V_low
+ 4.926000000e-07 V_low
+ 4.926010000e-07 V_low
+ 4.927000000e-07 V_low
+ 4.927010000e-07 V_low
+ 4.928000000e-07 V_low
+ 4.928010000e-07 V_low
+ 4.929000000e-07 V_low
+ 4.929010000e-07 V_hig
+ 4.930000000e-07 V_hig
+ 4.930010000e-07 V_hig
+ 4.931000000e-07 V_hig
+ 4.931010000e-07 V_hig
+ 4.932000000e-07 V_hig
+ 4.932010000e-07 V_hig
+ 4.933000000e-07 V_hig
+ 4.933010000e-07 V_hig
+ 4.934000000e-07 V_hig
+ 4.934010000e-07 V_hig
+ 4.935000000e-07 V_hig
+ 4.935010000e-07 V_hig
+ 4.936000000e-07 V_hig
+ 4.936010000e-07 V_hig
+ 4.937000000e-07 V_hig
+ 4.937010000e-07 V_hig
+ 4.938000000e-07 V_hig
+ 4.938010000e-07 V_hig
+ 4.939000000e-07 V_hig
+ 4.939010000e-07 V_hig
+ 4.940000000e-07 V_hig
+ 4.940010000e-07 V_hig
+ 4.941000000e-07 V_hig
+ 4.941010000e-07 V_hig
+ 4.942000000e-07 V_hig
+ 4.942010000e-07 V_hig
+ 4.943000000e-07 V_hig
+ 4.943010000e-07 V_hig
+ 4.944000000e-07 V_hig
+ 4.944010000e-07 V_hig
+ 4.945000000e-07 V_hig
+ 4.945010000e-07 V_hig
+ 4.946000000e-07 V_hig
+ 4.946010000e-07 V_hig
+ 4.947000000e-07 V_hig
+ 4.947010000e-07 V_hig
+ 4.948000000e-07 V_hig
+ 4.948010000e-07 V_hig
+ 4.949000000e-07 V_hig
+ 4.949010000e-07 V_low
+ 4.950000000e-07 V_low
+ 4.950010000e-07 V_low
+ 4.951000000e-07 V_low
+ 4.951010000e-07 V_low
+ 4.952000000e-07 V_low
+ 4.952010000e-07 V_low
+ 4.953000000e-07 V_low
+ 4.953010000e-07 V_low
+ 4.954000000e-07 V_low
+ 4.954010000e-07 V_low
+ 4.955000000e-07 V_low
+ 4.955010000e-07 V_low
+ 4.956000000e-07 V_low
+ 4.956010000e-07 V_low
+ 4.957000000e-07 V_low
+ 4.957010000e-07 V_low
+ 4.958000000e-07 V_low
+ 4.958010000e-07 V_low
+ 4.959000000e-07 V_low
+ 4.959010000e-07 V_low
+ 4.960000000e-07 V_low
+ 4.960010000e-07 V_low
+ 4.961000000e-07 V_low
+ 4.961010000e-07 V_low
+ 4.962000000e-07 V_low
+ 4.962010000e-07 V_low
+ 4.963000000e-07 V_low
+ 4.963010000e-07 V_low
+ 4.964000000e-07 V_low
+ 4.964010000e-07 V_low
+ 4.965000000e-07 V_low
+ 4.965010000e-07 V_low
+ 4.966000000e-07 V_low
+ 4.966010000e-07 V_low
+ 4.967000000e-07 V_low
+ 4.967010000e-07 V_low
+ 4.968000000e-07 V_low
+ 4.968010000e-07 V_low
+ 4.969000000e-07 V_low
+ 4.969010000e-07 V_hig
+ 4.970000000e-07 V_hig
+ 4.970010000e-07 V_hig
+ 4.971000000e-07 V_hig
+ 4.971010000e-07 V_hig
+ 4.972000000e-07 V_hig
+ 4.972010000e-07 V_hig
+ 4.973000000e-07 V_hig
+ 4.973010000e-07 V_hig
+ 4.974000000e-07 V_hig
+ 4.974010000e-07 V_hig
+ 4.975000000e-07 V_hig
+ 4.975010000e-07 V_hig
+ 4.976000000e-07 V_hig
+ 4.976010000e-07 V_hig
+ 4.977000000e-07 V_hig
+ 4.977010000e-07 V_hig
+ 4.978000000e-07 V_hig
+ 4.978010000e-07 V_hig
+ 4.979000000e-07 V_hig
+ 4.979010000e-07 V_hig
+ 4.980000000e-07 V_hig
+ 4.980010000e-07 V_hig
+ 4.981000000e-07 V_hig
+ 4.981010000e-07 V_hig
+ 4.982000000e-07 V_hig
+ 4.982010000e-07 V_hig
+ 4.983000000e-07 V_hig
+ 4.983010000e-07 V_hig
+ 4.984000000e-07 V_hig
+ 4.984010000e-07 V_hig
+ 4.985000000e-07 V_hig
+ 4.985010000e-07 V_hig
+ 4.986000000e-07 V_hig
+ 4.986010000e-07 V_hig
+ 4.987000000e-07 V_hig
+ 4.987010000e-07 V_hig
+ 4.988000000e-07 V_hig
+ 4.988010000e-07 V_hig
+ 4.989000000e-07 V_hig
+ 4.989010000e-07 V_hig
+ 4.990000000e-07 V_hig
+ 4.990010000e-07 V_hig
+ 4.991000000e-07 V_hig
+ 4.991010000e-07 V_hig
+ 4.992000000e-07 V_hig
+ 4.992010000e-07 V_hig
+ 4.993000000e-07 V_hig
+ 4.993010000e-07 V_hig
+ 4.994000000e-07 V_hig
+ 4.994010000e-07 V_hig
+ 4.995000000e-07 V_hig
+ 4.995010000e-07 V_hig
+ 4.996000000e-07 V_hig
+ 4.996010000e-07 V_hig
+ 4.997000000e-07 V_hig
+ 4.997010000e-07 V_hig
+ 4.998000000e-07 V_hig
+ 4.998010000e-07 V_hig
+ 4.999000000e-07 V_hig
+ 4.999010000e-07 V_low
+ 5.000000000e-07 V_low
+ 5.000010000e-07 V_low
+ 5.001000000e-07 V_low
+ 5.001010000e-07 V_low
+ 5.002000000e-07 V_low
+ 5.002010000e-07 V_low
+ 5.003000000e-07 V_low
+ 5.003010000e-07 V_low
+ 5.004000000e-07 V_low
+ 5.004010000e-07 V_low
+ 5.005000000e-07 V_low
+ 5.005010000e-07 V_low
+ 5.006000000e-07 V_low
+ 5.006010000e-07 V_low
+ 5.007000000e-07 V_low
+ 5.007010000e-07 V_low
+ 5.008000000e-07 V_low
+ 5.008010000e-07 V_low
+ 5.009000000e-07 V_low
+ 5.009010000e-07 V_hig
+ 5.010000000e-07 V_hig
+ 5.010010000e-07 V_hig
+ 5.011000000e-07 V_hig
+ 5.011010000e-07 V_hig
+ 5.012000000e-07 V_hig
+ 5.012010000e-07 V_hig
+ 5.013000000e-07 V_hig
+ 5.013010000e-07 V_hig
+ 5.014000000e-07 V_hig
+ 5.014010000e-07 V_hig
+ 5.015000000e-07 V_hig
+ 5.015010000e-07 V_hig
+ 5.016000000e-07 V_hig
+ 5.016010000e-07 V_hig
+ 5.017000000e-07 V_hig
+ 5.017010000e-07 V_hig
+ 5.018000000e-07 V_hig
+ 5.018010000e-07 V_hig
+ 5.019000000e-07 V_hig
+ 5.019010000e-07 V_hig
+ 5.020000000e-07 V_hig
+ 5.020010000e-07 V_hig
+ 5.021000000e-07 V_hig
+ 5.021010000e-07 V_hig
+ 5.022000000e-07 V_hig
+ 5.022010000e-07 V_hig
+ 5.023000000e-07 V_hig
+ 5.023010000e-07 V_hig
+ 5.024000000e-07 V_hig
+ 5.024010000e-07 V_hig
+ 5.025000000e-07 V_hig
+ 5.025010000e-07 V_hig
+ 5.026000000e-07 V_hig
+ 5.026010000e-07 V_hig
+ 5.027000000e-07 V_hig
+ 5.027010000e-07 V_hig
+ 5.028000000e-07 V_hig
+ 5.028010000e-07 V_hig
+ 5.029000000e-07 V_hig
+ 5.029010000e-07 V_hig
+ 5.030000000e-07 V_hig
+ 5.030010000e-07 V_hig
+ 5.031000000e-07 V_hig
+ 5.031010000e-07 V_hig
+ 5.032000000e-07 V_hig
+ 5.032010000e-07 V_hig
+ 5.033000000e-07 V_hig
+ 5.033010000e-07 V_hig
+ 5.034000000e-07 V_hig
+ 5.034010000e-07 V_hig
+ 5.035000000e-07 V_hig
+ 5.035010000e-07 V_hig
+ 5.036000000e-07 V_hig
+ 5.036010000e-07 V_hig
+ 5.037000000e-07 V_hig
+ 5.037010000e-07 V_hig
+ 5.038000000e-07 V_hig
+ 5.038010000e-07 V_hig
+ 5.039000000e-07 V_hig
+ 5.039010000e-07 V_low
+ 5.040000000e-07 V_low
+ 5.040010000e-07 V_low
+ 5.041000000e-07 V_low
+ 5.041010000e-07 V_low
+ 5.042000000e-07 V_low
+ 5.042010000e-07 V_low
+ 5.043000000e-07 V_low
+ 5.043010000e-07 V_low
+ 5.044000000e-07 V_low
+ 5.044010000e-07 V_low
+ 5.045000000e-07 V_low
+ 5.045010000e-07 V_low
+ 5.046000000e-07 V_low
+ 5.046010000e-07 V_low
+ 5.047000000e-07 V_low
+ 5.047010000e-07 V_low
+ 5.048000000e-07 V_low
+ 5.048010000e-07 V_low
+ 5.049000000e-07 V_low
+ 5.049010000e-07 V_low
+ 5.050000000e-07 V_low
+ 5.050010000e-07 V_low
+ 5.051000000e-07 V_low
+ 5.051010000e-07 V_low
+ 5.052000000e-07 V_low
+ 5.052010000e-07 V_low
+ 5.053000000e-07 V_low
+ 5.053010000e-07 V_low
+ 5.054000000e-07 V_low
+ 5.054010000e-07 V_low
+ 5.055000000e-07 V_low
+ 5.055010000e-07 V_low
+ 5.056000000e-07 V_low
+ 5.056010000e-07 V_low
+ 5.057000000e-07 V_low
+ 5.057010000e-07 V_low
+ 5.058000000e-07 V_low
+ 5.058010000e-07 V_low
+ 5.059000000e-07 V_low
+ 5.059010000e-07 V_low
+ 5.060000000e-07 V_low
+ 5.060010000e-07 V_low
+ 5.061000000e-07 V_low
+ 5.061010000e-07 V_low
+ 5.062000000e-07 V_low
+ 5.062010000e-07 V_low
+ 5.063000000e-07 V_low
+ 5.063010000e-07 V_low
+ 5.064000000e-07 V_low
+ 5.064010000e-07 V_low
+ 5.065000000e-07 V_low
+ 5.065010000e-07 V_low
+ 5.066000000e-07 V_low
+ 5.066010000e-07 V_low
+ 5.067000000e-07 V_low
+ 5.067010000e-07 V_low
+ 5.068000000e-07 V_low
+ 5.068010000e-07 V_low
+ 5.069000000e-07 V_low
+ 5.069010000e-07 V_hig
+ 5.070000000e-07 V_hig
+ 5.070010000e-07 V_hig
+ 5.071000000e-07 V_hig
+ 5.071010000e-07 V_hig
+ 5.072000000e-07 V_hig
+ 5.072010000e-07 V_hig
+ 5.073000000e-07 V_hig
+ 5.073010000e-07 V_hig
+ 5.074000000e-07 V_hig
+ 5.074010000e-07 V_hig
+ 5.075000000e-07 V_hig
+ 5.075010000e-07 V_hig
+ 5.076000000e-07 V_hig
+ 5.076010000e-07 V_hig
+ 5.077000000e-07 V_hig
+ 5.077010000e-07 V_hig
+ 5.078000000e-07 V_hig
+ 5.078010000e-07 V_hig
+ 5.079000000e-07 V_hig
+ 5.079010000e-07 V_hig
+ 5.080000000e-07 V_hig
+ 5.080010000e-07 V_hig
+ 5.081000000e-07 V_hig
+ 5.081010000e-07 V_hig
+ 5.082000000e-07 V_hig
+ 5.082010000e-07 V_hig
+ 5.083000000e-07 V_hig
+ 5.083010000e-07 V_hig
+ 5.084000000e-07 V_hig
+ 5.084010000e-07 V_hig
+ 5.085000000e-07 V_hig
+ 5.085010000e-07 V_hig
+ 5.086000000e-07 V_hig
+ 5.086010000e-07 V_hig
+ 5.087000000e-07 V_hig
+ 5.087010000e-07 V_hig
+ 5.088000000e-07 V_hig
+ 5.088010000e-07 V_hig
+ 5.089000000e-07 V_hig
+ 5.089010000e-07 V_hig
+ 5.090000000e-07 V_hig
+ 5.090010000e-07 V_hig
+ 5.091000000e-07 V_hig
+ 5.091010000e-07 V_hig
+ 5.092000000e-07 V_hig
+ 5.092010000e-07 V_hig
+ 5.093000000e-07 V_hig
+ 5.093010000e-07 V_hig
+ 5.094000000e-07 V_hig
+ 5.094010000e-07 V_hig
+ 5.095000000e-07 V_hig
+ 5.095010000e-07 V_hig
+ 5.096000000e-07 V_hig
+ 5.096010000e-07 V_hig
+ 5.097000000e-07 V_hig
+ 5.097010000e-07 V_hig
+ 5.098000000e-07 V_hig
+ 5.098010000e-07 V_hig
+ 5.099000000e-07 V_hig
+ 5.099010000e-07 V_low
+ 5.100000000e-07 V_low
+ 5.100010000e-07 V_low
+ 5.101000000e-07 V_low
+ 5.101010000e-07 V_low
+ 5.102000000e-07 V_low
+ 5.102010000e-07 V_low
+ 5.103000000e-07 V_low
+ 5.103010000e-07 V_low
+ 5.104000000e-07 V_low
+ 5.104010000e-07 V_low
+ 5.105000000e-07 V_low
+ 5.105010000e-07 V_low
+ 5.106000000e-07 V_low
+ 5.106010000e-07 V_low
+ 5.107000000e-07 V_low
+ 5.107010000e-07 V_low
+ 5.108000000e-07 V_low
+ 5.108010000e-07 V_low
+ 5.109000000e-07 V_low
+ 5.109010000e-07 V_low
+ 5.110000000e-07 V_low
+ 5.110010000e-07 V_low
+ 5.111000000e-07 V_low
+ 5.111010000e-07 V_low
+ 5.112000000e-07 V_low
+ 5.112010000e-07 V_low
+ 5.113000000e-07 V_low
+ 5.113010000e-07 V_low
+ 5.114000000e-07 V_low
+ 5.114010000e-07 V_low
+ 5.115000000e-07 V_low
+ 5.115010000e-07 V_low
+ 5.116000000e-07 V_low
+ 5.116010000e-07 V_low
+ 5.117000000e-07 V_low
+ 5.117010000e-07 V_low
+ 5.118000000e-07 V_low
+ 5.118010000e-07 V_low
+ 5.119000000e-07 V_low
+ 5.119010000e-07 V_low
+ 5.120000000e-07 V_low
+ 5.120010000e-07 V_low
+ 5.121000000e-07 V_low
+ 5.121010000e-07 V_low
+ 5.122000000e-07 V_low
+ 5.122010000e-07 V_low
+ 5.123000000e-07 V_low
+ 5.123010000e-07 V_low
+ 5.124000000e-07 V_low
+ 5.124010000e-07 V_low
+ 5.125000000e-07 V_low
+ 5.125010000e-07 V_low
+ 5.126000000e-07 V_low
+ 5.126010000e-07 V_low
+ 5.127000000e-07 V_low
+ 5.127010000e-07 V_low
+ 5.128000000e-07 V_low
+ 5.128010000e-07 V_low
+ 5.129000000e-07 V_low
+ 5.129010000e-07 V_hig
+ 5.130000000e-07 V_hig
+ 5.130010000e-07 V_hig
+ 5.131000000e-07 V_hig
+ 5.131010000e-07 V_hig
+ 5.132000000e-07 V_hig
+ 5.132010000e-07 V_hig
+ 5.133000000e-07 V_hig
+ 5.133010000e-07 V_hig
+ 5.134000000e-07 V_hig
+ 5.134010000e-07 V_hig
+ 5.135000000e-07 V_hig
+ 5.135010000e-07 V_hig
+ 5.136000000e-07 V_hig
+ 5.136010000e-07 V_hig
+ 5.137000000e-07 V_hig
+ 5.137010000e-07 V_hig
+ 5.138000000e-07 V_hig
+ 5.138010000e-07 V_hig
+ 5.139000000e-07 V_hig
+ 5.139010000e-07 V_hig
+ 5.140000000e-07 V_hig
+ 5.140010000e-07 V_hig
+ 5.141000000e-07 V_hig
+ 5.141010000e-07 V_hig
+ 5.142000000e-07 V_hig
+ 5.142010000e-07 V_hig
+ 5.143000000e-07 V_hig
+ 5.143010000e-07 V_hig
+ 5.144000000e-07 V_hig
+ 5.144010000e-07 V_hig
+ 5.145000000e-07 V_hig
+ 5.145010000e-07 V_hig
+ 5.146000000e-07 V_hig
+ 5.146010000e-07 V_hig
+ 5.147000000e-07 V_hig
+ 5.147010000e-07 V_hig
+ 5.148000000e-07 V_hig
+ 5.148010000e-07 V_hig
+ 5.149000000e-07 V_hig
+ 5.149010000e-07 V_low
+ 5.150000000e-07 V_low
+ 5.150010000e-07 V_low
+ 5.151000000e-07 V_low
+ 5.151010000e-07 V_low
+ 5.152000000e-07 V_low
+ 5.152010000e-07 V_low
+ 5.153000000e-07 V_low
+ 5.153010000e-07 V_low
+ 5.154000000e-07 V_low
+ 5.154010000e-07 V_low
+ 5.155000000e-07 V_low
+ 5.155010000e-07 V_low
+ 5.156000000e-07 V_low
+ 5.156010000e-07 V_low
+ 5.157000000e-07 V_low
+ 5.157010000e-07 V_low
+ 5.158000000e-07 V_low
+ 5.158010000e-07 V_low
+ 5.159000000e-07 V_low
+ 5.159010000e-07 V_low
+ 5.160000000e-07 V_low
+ 5.160010000e-07 V_low
+ 5.161000000e-07 V_low
+ 5.161010000e-07 V_low
+ 5.162000000e-07 V_low
+ 5.162010000e-07 V_low
+ 5.163000000e-07 V_low
+ 5.163010000e-07 V_low
+ 5.164000000e-07 V_low
+ 5.164010000e-07 V_low
+ 5.165000000e-07 V_low
+ 5.165010000e-07 V_low
+ 5.166000000e-07 V_low
+ 5.166010000e-07 V_low
+ 5.167000000e-07 V_low
+ 5.167010000e-07 V_low
+ 5.168000000e-07 V_low
+ 5.168010000e-07 V_low
+ 5.169000000e-07 V_low
+ 5.169010000e-07 V_hig
+ 5.170000000e-07 V_hig
+ 5.170010000e-07 V_hig
+ 5.171000000e-07 V_hig
+ 5.171010000e-07 V_hig
+ 5.172000000e-07 V_hig
+ 5.172010000e-07 V_hig
+ 5.173000000e-07 V_hig
+ 5.173010000e-07 V_hig
+ 5.174000000e-07 V_hig
+ 5.174010000e-07 V_hig
+ 5.175000000e-07 V_hig
+ 5.175010000e-07 V_hig
+ 5.176000000e-07 V_hig
+ 5.176010000e-07 V_hig
+ 5.177000000e-07 V_hig
+ 5.177010000e-07 V_hig
+ 5.178000000e-07 V_hig
+ 5.178010000e-07 V_hig
+ 5.179000000e-07 V_hig
+ 5.179010000e-07 V_hig
+ 5.180000000e-07 V_hig
+ 5.180010000e-07 V_hig
+ 5.181000000e-07 V_hig
+ 5.181010000e-07 V_hig
+ 5.182000000e-07 V_hig
+ 5.182010000e-07 V_hig
+ 5.183000000e-07 V_hig
+ 5.183010000e-07 V_hig
+ 5.184000000e-07 V_hig
+ 5.184010000e-07 V_hig
+ 5.185000000e-07 V_hig
+ 5.185010000e-07 V_hig
+ 5.186000000e-07 V_hig
+ 5.186010000e-07 V_hig
+ 5.187000000e-07 V_hig
+ 5.187010000e-07 V_hig
+ 5.188000000e-07 V_hig
+ 5.188010000e-07 V_hig
+ 5.189000000e-07 V_hig
+ 5.189010000e-07 V_hig
+ 5.190000000e-07 V_hig
+ 5.190010000e-07 V_hig
+ 5.191000000e-07 V_hig
+ 5.191010000e-07 V_hig
+ 5.192000000e-07 V_hig
+ 5.192010000e-07 V_hig
+ 5.193000000e-07 V_hig
+ 5.193010000e-07 V_hig
+ 5.194000000e-07 V_hig
+ 5.194010000e-07 V_hig
+ 5.195000000e-07 V_hig
+ 5.195010000e-07 V_hig
+ 5.196000000e-07 V_hig
+ 5.196010000e-07 V_hig
+ 5.197000000e-07 V_hig
+ 5.197010000e-07 V_hig
+ 5.198000000e-07 V_hig
+ 5.198010000e-07 V_hig
+ 5.199000000e-07 V_hig
+ 5.199010000e-07 V_hig
+ 5.200000000e-07 V_hig
+ 5.200010000e-07 V_hig
+ 5.201000000e-07 V_hig
+ 5.201010000e-07 V_hig
+ 5.202000000e-07 V_hig
+ 5.202010000e-07 V_hig
+ 5.203000000e-07 V_hig
+ 5.203010000e-07 V_hig
+ 5.204000000e-07 V_hig
+ 5.204010000e-07 V_hig
+ 5.205000000e-07 V_hig
+ 5.205010000e-07 V_hig
+ 5.206000000e-07 V_hig
+ 5.206010000e-07 V_hig
+ 5.207000000e-07 V_hig
+ 5.207010000e-07 V_hig
+ 5.208000000e-07 V_hig
+ 5.208010000e-07 V_hig
+ 5.209000000e-07 V_hig
+ 5.209010000e-07 V_hig
+ 5.210000000e-07 V_hig
+ 5.210010000e-07 V_hig
+ 5.211000000e-07 V_hig
+ 5.211010000e-07 V_hig
+ 5.212000000e-07 V_hig
+ 5.212010000e-07 V_hig
+ 5.213000000e-07 V_hig
+ 5.213010000e-07 V_hig
+ 5.214000000e-07 V_hig
+ 5.214010000e-07 V_hig
+ 5.215000000e-07 V_hig
+ 5.215010000e-07 V_hig
+ 5.216000000e-07 V_hig
+ 5.216010000e-07 V_hig
+ 5.217000000e-07 V_hig
+ 5.217010000e-07 V_hig
+ 5.218000000e-07 V_hig
+ 5.218010000e-07 V_hig
+ 5.219000000e-07 V_hig
+ 5.219010000e-07 V_hig
+ 5.220000000e-07 V_hig
+ 5.220010000e-07 V_hig
+ 5.221000000e-07 V_hig
+ 5.221010000e-07 V_hig
+ 5.222000000e-07 V_hig
+ 5.222010000e-07 V_hig
+ 5.223000000e-07 V_hig
+ 5.223010000e-07 V_hig
+ 5.224000000e-07 V_hig
+ 5.224010000e-07 V_hig
+ 5.225000000e-07 V_hig
+ 5.225010000e-07 V_hig
+ 5.226000000e-07 V_hig
+ 5.226010000e-07 V_hig
+ 5.227000000e-07 V_hig
+ 5.227010000e-07 V_hig
+ 5.228000000e-07 V_hig
+ 5.228010000e-07 V_hig
+ 5.229000000e-07 V_hig
+ 5.229010000e-07 V_low
+ 5.230000000e-07 V_low
+ 5.230010000e-07 V_low
+ 5.231000000e-07 V_low
+ 5.231010000e-07 V_low
+ 5.232000000e-07 V_low
+ 5.232010000e-07 V_low
+ 5.233000000e-07 V_low
+ 5.233010000e-07 V_low
+ 5.234000000e-07 V_low
+ 5.234010000e-07 V_low
+ 5.235000000e-07 V_low
+ 5.235010000e-07 V_low
+ 5.236000000e-07 V_low
+ 5.236010000e-07 V_low
+ 5.237000000e-07 V_low
+ 5.237010000e-07 V_low
+ 5.238000000e-07 V_low
+ 5.238010000e-07 V_low
+ 5.239000000e-07 V_low
+ 5.239010000e-07 V_low
+ 5.240000000e-07 V_low
+ 5.240010000e-07 V_low
+ 5.241000000e-07 V_low
+ 5.241010000e-07 V_low
+ 5.242000000e-07 V_low
+ 5.242010000e-07 V_low
+ 5.243000000e-07 V_low
+ 5.243010000e-07 V_low
+ 5.244000000e-07 V_low
+ 5.244010000e-07 V_low
+ 5.245000000e-07 V_low
+ 5.245010000e-07 V_low
+ 5.246000000e-07 V_low
+ 5.246010000e-07 V_low
+ 5.247000000e-07 V_low
+ 5.247010000e-07 V_low
+ 5.248000000e-07 V_low
+ 5.248010000e-07 V_low
+ 5.249000000e-07 V_low
+ 5.249010000e-07 V_low
+ 5.250000000e-07 V_low
+ 5.250010000e-07 V_low
+ 5.251000000e-07 V_low
+ 5.251010000e-07 V_low
+ 5.252000000e-07 V_low
+ 5.252010000e-07 V_low
+ 5.253000000e-07 V_low
+ 5.253010000e-07 V_low
+ 5.254000000e-07 V_low
+ 5.254010000e-07 V_low
+ 5.255000000e-07 V_low
+ 5.255010000e-07 V_low
+ 5.256000000e-07 V_low
+ 5.256010000e-07 V_low
+ 5.257000000e-07 V_low
+ 5.257010000e-07 V_low
+ 5.258000000e-07 V_low
+ 5.258010000e-07 V_low
+ 5.259000000e-07 V_low
+ 5.259010000e-07 V_hig
+ 5.260000000e-07 V_hig
+ 5.260010000e-07 V_hig
+ 5.261000000e-07 V_hig
+ 5.261010000e-07 V_hig
+ 5.262000000e-07 V_hig
+ 5.262010000e-07 V_hig
+ 5.263000000e-07 V_hig
+ 5.263010000e-07 V_hig
+ 5.264000000e-07 V_hig
+ 5.264010000e-07 V_hig
+ 5.265000000e-07 V_hig
+ 5.265010000e-07 V_hig
+ 5.266000000e-07 V_hig
+ 5.266010000e-07 V_hig
+ 5.267000000e-07 V_hig
+ 5.267010000e-07 V_hig
+ 5.268000000e-07 V_hig
+ 5.268010000e-07 V_hig
+ 5.269000000e-07 V_hig
+ 5.269010000e-07 V_low
+ 5.270000000e-07 V_low
+ 5.270010000e-07 V_low
+ 5.271000000e-07 V_low
+ 5.271010000e-07 V_low
+ 5.272000000e-07 V_low
+ 5.272010000e-07 V_low
+ 5.273000000e-07 V_low
+ 5.273010000e-07 V_low
+ 5.274000000e-07 V_low
+ 5.274010000e-07 V_low
+ 5.275000000e-07 V_low
+ 5.275010000e-07 V_low
+ 5.276000000e-07 V_low
+ 5.276010000e-07 V_low
+ 5.277000000e-07 V_low
+ 5.277010000e-07 V_low
+ 5.278000000e-07 V_low
+ 5.278010000e-07 V_low
+ 5.279000000e-07 V_low
+ 5.279010000e-07 V_low
+ 5.280000000e-07 V_low
+ 5.280010000e-07 V_low
+ 5.281000000e-07 V_low
+ 5.281010000e-07 V_low
+ 5.282000000e-07 V_low
+ 5.282010000e-07 V_low
+ 5.283000000e-07 V_low
+ 5.283010000e-07 V_low
+ 5.284000000e-07 V_low
+ 5.284010000e-07 V_low
+ 5.285000000e-07 V_low
+ 5.285010000e-07 V_low
+ 5.286000000e-07 V_low
+ 5.286010000e-07 V_low
+ 5.287000000e-07 V_low
+ 5.287010000e-07 V_low
+ 5.288000000e-07 V_low
+ 5.288010000e-07 V_low
+ 5.289000000e-07 V_low
+ 5.289010000e-07 V_low
+ 5.290000000e-07 V_low
+ 5.290010000e-07 V_low
+ 5.291000000e-07 V_low
+ 5.291010000e-07 V_low
+ 5.292000000e-07 V_low
+ 5.292010000e-07 V_low
+ 5.293000000e-07 V_low
+ 5.293010000e-07 V_low
+ 5.294000000e-07 V_low
+ 5.294010000e-07 V_low
+ 5.295000000e-07 V_low
+ 5.295010000e-07 V_low
+ 5.296000000e-07 V_low
+ 5.296010000e-07 V_low
+ 5.297000000e-07 V_low
+ 5.297010000e-07 V_low
+ 5.298000000e-07 V_low
+ 5.298010000e-07 V_low
+ 5.299000000e-07 V_low
+ 5.299010000e-07 V_hig
+ 5.300000000e-07 V_hig
+ 5.300010000e-07 V_hig
+ 5.301000000e-07 V_hig
+ 5.301010000e-07 V_hig
+ 5.302000000e-07 V_hig
+ 5.302010000e-07 V_hig
+ 5.303000000e-07 V_hig
+ 5.303010000e-07 V_hig
+ 5.304000000e-07 V_hig
+ 5.304010000e-07 V_hig
+ 5.305000000e-07 V_hig
+ 5.305010000e-07 V_hig
+ 5.306000000e-07 V_hig
+ 5.306010000e-07 V_hig
+ 5.307000000e-07 V_hig
+ 5.307010000e-07 V_hig
+ 5.308000000e-07 V_hig
+ 5.308010000e-07 V_hig
+ 5.309000000e-07 V_hig
+ 5.309010000e-07 V_hig
+ 5.310000000e-07 V_hig
+ 5.310010000e-07 V_hig
+ 5.311000000e-07 V_hig
+ 5.311010000e-07 V_hig
+ 5.312000000e-07 V_hig
+ 5.312010000e-07 V_hig
+ 5.313000000e-07 V_hig
+ 5.313010000e-07 V_hig
+ 5.314000000e-07 V_hig
+ 5.314010000e-07 V_hig
+ 5.315000000e-07 V_hig
+ 5.315010000e-07 V_hig
+ 5.316000000e-07 V_hig
+ 5.316010000e-07 V_hig
+ 5.317000000e-07 V_hig
+ 5.317010000e-07 V_hig
+ 5.318000000e-07 V_hig
+ 5.318010000e-07 V_hig
+ 5.319000000e-07 V_hig
+ 5.319010000e-07 V_hig
+ 5.320000000e-07 V_hig
+ 5.320010000e-07 V_hig
+ 5.321000000e-07 V_hig
+ 5.321010000e-07 V_hig
+ 5.322000000e-07 V_hig
+ 5.322010000e-07 V_hig
+ 5.323000000e-07 V_hig
+ 5.323010000e-07 V_hig
+ 5.324000000e-07 V_hig
+ 5.324010000e-07 V_hig
+ 5.325000000e-07 V_hig
+ 5.325010000e-07 V_hig
+ 5.326000000e-07 V_hig
+ 5.326010000e-07 V_hig
+ 5.327000000e-07 V_hig
+ 5.327010000e-07 V_hig
+ 5.328000000e-07 V_hig
+ 5.328010000e-07 V_hig
+ 5.329000000e-07 V_hig
+ 5.329010000e-07 V_low
+ 5.330000000e-07 V_low
+ 5.330010000e-07 V_low
+ 5.331000000e-07 V_low
+ 5.331010000e-07 V_low
+ 5.332000000e-07 V_low
+ 5.332010000e-07 V_low
+ 5.333000000e-07 V_low
+ 5.333010000e-07 V_low
+ 5.334000000e-07 V_low
+ 5.334010000e-07 V_low
+ 5.335000000e-07 V_low
+ 5.335010000e-07 V_low
+ 5.336000000e-07 V_low
+ 5.336010000e-07 V_low
+ 5.337000000e-07 V_low
+ 5.337010000e-07 V_low
+ 5.338000000e-07 V_low
+ 5.338010000e-07 V_low
+ 5.339000000e-07 V_low
+ 5.339010000e-07 V_hig
+ 5.340000000e-07 V_hig
+ 5.340010000e-07 V_hig
+ 5.341000000e-07 V_hig
+ 5.341010000e-07 V_hig
+ 5.342000000e-07 V_hig
+ 5.342010000e-07 V_hig
+ 5.343000000e-07 V_hig
+ 5.343010000e-07 V_hig
+ 5.344000000e-07 V_hig
+ 5.344010000e-07 V_hig
+ 5.345000000e-07 V_hig
+ 5.345010000e-07 V_hig
+ 5.346000000e-07 V_hig
+ 5.346010000e-07 V_hig
+ 5.347000000e-07 V_hig
+ 5.347010000e-07 V_hig
+ 5.348000000e-07 V_hig
+ 5.348010000e-07 V_hig
+ 5.349000000e-07 V_hig
+ 5.349010000e-07 V_hig
+ 5.350000000e-07 V_hig
+ 5.350010000e-07 V_hig
+ 5.351000000e-07 V_hig
+ 5.351010000e-07 V_hig
+ 5.352000000e-07 V_hig
+ 5.352010000e-07 V_hig
+ 5.353000000e-07 V_hig
+ 5.353010000e-07 V_hig
+ 5.354000000e-07 V_hig
+ 5.354010000e-07 V_hig
+ 5.355000000e-07 V_hig
+ 5.355010000e-07 V_hig
+ 5.356000000e-07 V_hig
+ 5.356010000e-07 V_hig
+ 5.357000000e-07 V_hig
+ 5.357010000e-07 V_hig
+ 5.358000000e-07 V_hig
+ 5.358010000e-07 V_hig
+ 5.359000000e-07 V_hig
+ 5.359010000e-07 V_hig
+ 5.360000000e-07 V_hig
+ 5.360010000e-07 V_hig
+ 5.361000000e-07 V_hig
+ 5.361010000e-07 V_hig
+ 5.362000000e-07 V_hig
+ 5.362010000e-07 V_hig
+ 5.363000000e-07 V_hig
+ 5.363010000e-07 V_hig
+ 5.364000000e-07 V_hig
+ 5.364010000e-07 V_hig
+ 5.365000000e-07 V_hig
+ 5.365010000e-07 V_hig
+ 5.366000000e-07 V_hig
+ 5.366010000e-07 V_hig
+ 5.367000000e-07 V_hig
+ 5.367010000e-07 V_hig
+ 5.368000000e-07 V_hig
+ 5.368010000e-07 V_hig
+ 5.369000000e-07 V_hig
+ 5.369010000e-07 V_low
+ 5.370000000e-07 V_low
+ 5.370010000e-07 V_low
+ 5.371000000e-07 V_low
+ 5.371010000e-07 V_low
+ 5.372000000e-07 V_low
+ 5.372010000e-07 V_low
+ 5.373000000e-07 V_low
+ 5.373010000e-07 V_low
+ 5.374000000e-07 V_low
+ 5.374010000e-07 V_low
+ 5.375000000e-07 V_low
+ 5.375010000e-07 V_low
+ 5.376000000e-07 V_low
+ 5.376010000e-07 V_low
+ 5.377000000e-07 V_low
+ 5.377010000e-07 V_low
+ 5.378000000e-07 V_low
+ 5.378010000e-07 V_low
+ 5.379000000e-07 V_low
+ 5.379010000e-07 V_low
+ 5.380000000e-07 V_low
+ 5.380010000e-07 V_low
+ 5.381000000e-07 V_low
+ 5.381010000e-07 V_low
+ 5.382000000e-07 V_low
+ 5.382010000e-07 V_low
+ 5.383000000e-07 V_low
+ 5.383010000e-07 V_low
+ 5.384000000e-07 V_low
+ 5.384010000e-07 V_low
+ 5.385000000e-07 V_low
+ 5.385010000e-07 V_low
+ 5.386000000e-07 V_low
+ 5.386010000e-07 V_low
+ 5.387000000e-07 V_low
+ 5.387010000e-07 V_low
+ 5.388000000e-07 V_low
+ 5.388010000e-07 V_low
+ 5.389000000e-07 V_low
+ 5.389010000e-07 V_low
+ 5.390000000e-07 V_low
+ 5.390010000e-07 V_low
+ 5.391000000e-07 V_low
+ 5.391010000e-07 V_low
+ 5.392000000e-07 V_low
+ 5.392010000e-07 V_low
+ 5.393000000e-07 V_low
+ 5.393010000e-07 V_low
+ 5.394000000e-07 V_low
+ 5.394010000e-07 V_low
+ 5.395000000e-07 V_low
+ 5.395010000e-07 V_low
+ 5.396000000e-07 V_low
+ 5.396010000e-07 V_low
+ 5.397000000e-07 V_low
+ 5.397010000e-07 V_low
+ 5.398000000e-07 V_low
+ 5.398010000e-07 V_low
+ 5.399000000e-07 V_low
+ 5.399010000e-07 V_hig
+ 5.400000000e-07 V_hig
+ 5.400010000e-07 V_hig
+ 5.401000000e-07 V_hig
+ 5.401010000e-07 V_hig
+ 5.402000000e-07 V_hig
+ 5.402010000e-07 V_hig
+ 5.403000000e-07 V_hig
+ 5.403010000e-07 V_hig
+ 5.404000000e-07 V_hig
+ 5.404010000e-07 V_hig
+ 5.405000000e-07 V_hig
+ 5.405010000e-07 V_hig
+ 5.406000000e-07 V_hig
+ 5.406010000e-07 V_hig
+ 5.407000000e-07 V_hig
+ 5.407010000e-07 V_hig
+ 5.408000000e-07 V_hig
+ 5.408010000e-07 V_hig
+ 5.409000000e-07 V_hig
+ 5.409010000e-07 V_hig
+ 5.410000000e-07 V_hig
+ 5.410010000e-07 V_hig
+ 5.411000000e-07 V_hig
+ 5.411010000e-07 V_hig
+ 5.412000000e-07 V_hig
+ 5.412010000e-07 V_hig
+ 5.413000000e-07 V_hig
+ 5.413010000e-07 V_hig
+ 5.414000000e-07 V_hig
+ 5.414010000e-07 V_hig
+ 5.415000000e-07 V_hig
+ 5.415010000e-07 V_hig
+ 5.416000000e-07 V_hig
+ 5.416010000e-07 V_hig
+ 5.417000000e-07 V_hig
+ 5.417010000e-07 V_hig
+ 5.418000000e-07 V_hig
+ 5.418010000e-07 V_hig
+ 5.419000000e-07 V_hig
+ 5.419010000e-07 V_hig
+ 5.420000000e-07 V_hig
+ 5.420010000e-07 V_hig
+ 5.421000000e-07 V_hig
+ 5.421010000e-07 V_hig
+ 5.422000000e-07 V_hig
+ 5.422010000e-07 V_hig
+ 5.423000000e-07 V_hig
+ 5.423010000e-07 V_hig
+ 5.424000000e-07 V_hig
+ 5.424010000e-07 V_hig
+ 5.425000000e-07 V_hig
+ 5.425010000e-07 V_hig
+ 5.426000000e-07 V_hig
+ 5.426010000e-07 V_hig
+ 5.427000000e-07 V_hig
+ 5.427010000e-07 V_hig
+ 5.428000000e-07 V_hig
+ 5.428010000e-07 V_hig
+ 5.429000000e-07 V_hig
+ 5.429010000e-07 V_hig
+ 5.430000000e-07 V_hig
+ 5.430010000e-07 V_hig
+ 5.431000000e-07 V_hig
+ 5.431010000e-07 V_hig
+ 5.432000000e-07 V_hig
+ 5.432010000e-07 V_hig
+ 5.433000000e-07 V_hig
+ 5.433010000e-07 V_hig
+ 5.434000000e-07 V_hig
+ 5.434010000e-07 V_hig
+ 5.435000000e-07 V_hig
+ 5.435010000e-07 V_hig
+ 5.436000000e-07 V_hig
+ 5.436010000e-07 V_hig
+ 5.437000000e-07 V_hig
+ 5.437010000e-07 V_hig
+ 5.438000000e-07 V_hig
+ 5.438010000e-07 V_hig
+ 5.439000000e-07 V_hig
+ 5.439010000e-07 V_low
+ 5.440000000e-07 V_low
+ 5.440010000e-07 V_low
+ 5.441000000e-07 V_low
+ 5.441010000e-07 V_low
+ 5.442000000e-07 V_low
+ 5.442010000e-07 V_low
+ 5.443000000e-07 V_low
+ 5.443010000e-07 V_low
+ 5.444000000e-07 V_low
+ 5.444010000e-07 V_low
+ 5.445000000e-07 V_low
+ 5.445010000e-07 V_low
+ 5.446000000e-07 V_low
+ 5.446010000e-07 V_low
+ 5.447000000e-07 V_low
+ 5.447010000e-07 V_low
+ 5.448000000e-07 V_low
+ 5.448010000e-07 V_low
+ 5.449000000e-07 V_low
+ 5.449010000e-07 V_hig
+ 5.450000000e-07 V_hig
+ 5.450010000e-07 V_hig
+ 5.451000000e-07 V_hig
+ 5.451010000e-07 V_hig
+ 5.452000000e-07 V_hig
+ 5.452010000e-07 V_hig
+ 5.453000000e-07 V_hig
+ 5.453010000e-07 V_hig
+ 5.454000000e-07 V_hig
+ 5.454010000e-07 V_hig
+ 5.455000000e-07 V_hig
+ 5.455010000e-07 V_hig
+ 5.456000000e-07 V_hig
+ 5.456010000e-07 V_hig
+ 5.457000000e-07 V_hig
+ 5.457010000e-07 V_hig
+ 5.458000000e-07 V_hig
+ 5.458010000e-07 V_hig
+ 5.459000000e-07 V_hig
+ 5.459010000e-07 V_hig
+ 5.460000000e-07 V_hig
+ 5.460010000e-07 V_hig
+ 5.461000000e-07 V_hig
+ 5.461010000e-07 V_hig
+ 5.462000000e-07 V_hig
+ 5.462010000e-07 V_hig
+ 5.463000000e-07 V_hig
+ 5.463010000e-07 V_hig
+ 5.464000000e-07 V_hig
+ 5.464010000e-07 V_hig
+ 5.465000000e-07 V_hig
+ 5.465010000e-07 V_hig
+ 5.466000000e-07 V_hig
+ 5.466010000e-07 V_hig
+ 5.467000000e-07 V_hig
+ 5.467010000e-07 V_hig
+ 5.468000000e-07 V_hig
+ 5.468010000e-07 V_hig
+ 5.469000000e-07 V_hig
+ 5.469010000e-07 V_hig
+ 5.470000000e-07 V_hig
+ 5.470010000e-07 V_hig
+ 5.471000000e-07 V_hig
+ 5.471010000e-07 V_hig
+ 5.472000000e-07 V_hig
+ 5.472010000e-07 V_hig
+ 5.473000000e-07 V_hig
+ 5.473010000e-07 V_hig
+ 5.474000000e-07 V_hig
+ 5.474010000e-07 V_hig
+ 5.475000000e-07 V_hig
+ 5.475010000e-07 V_hig
+ 5.476000000e-07 V_hig
+ 5.476010000e-07 V_hig
+ 5.477000000e-07 V_hig
+ 5.477010000e-07 V_hig
+ 5.478000000e-07 V_hig
+ 5.478010000e-07 V_hig
+ 5.479000000e-07 V_hig
+ 5.479010000e-07 V_low
+ 5.480000000e-07 V_low
+ 5.480010000e-07 V_low
+ 5.481000000e-07 V_low
+ 5.481010000e-07 V_low
+ 5.482000000e-07 V_low
+ 5.482010000e-07 V_low
+ 5.483000000e-07 V_low
+ 5.483010000e-07 V_low
+ 5.484000000e-07 V_low
+ 5.484010000e-07 V_low
+ 5.485000000e-07 V_low
+ 5.485010000e-07 V_low
+ 5.486000000e-07 V_low
+ 5.486010000e-07 V_low
+ 5.487000000e-07 V_low
+ 5.487010000e-07 V_low
+ 5.488000000e-07 V_low
+ 5.488010000e-07 V_low
+ 5.489000000e-07 V_low
+ 5.489010000e-07 V_hig
+ 5.490000000e-07 V_hig
+ 5.490010000e-07 V_hig
+ 5.491000000e-07 V_hig
+ 5.491010000e-07 V_hig
+ 5.492000000e-07 V_hig
+ 5.492010000e-07 V_hig
+ 5.493000000e-07 V_hig
+ 5.493010000e-07 V_hig
+ 5.494000000e-07 V_hig
+ 5.494010000e-07 V_hig
+ 5.495000000e-07 V_hig
+ 5.495010000e-07 V_hig
+ 5.496000000e-07 V_hig
+ 5.496010000e-07 V_hig
+ 5.497000000e-07 V_hig
+ 5.497010000e-07 V_hig
+ 5.498000000e-07 V_hig
+ 5.498010000e-07 V_hig
+ 5.499000000e-07 V_hig
+ 5.499010000e-07 V_hig
+ 5.500000000e-07 V_hig
+ 5.500010000e-07 V_hig
+ 5.501000000e-07 V_hig
+ 5.501010000e-07 V_hig
+ 5.502000000e-07 V_hig
+ 5.502010000e-07 V_hig
+ 5.503000000e-07 V_hig
+ 5.503010000e-07 V_hig
+ 5.504000000e-07 V_hig
+ 5.504010000e-07 V_hig
+ 5.505000000e-07 V_hig
+ 5.505010000e-07 V_hig
+ 5.506000000e-07 V_hig
+ 5.506010000e-07 V_hig
+ 5.507000000e-07 V_hig
+ 5.507010000e-07 V_hig
+ 5.508000000e-07 V_hig
+ 5.508010000e-07 V_hig
+ 5.509000000e-07 V_hig
+ 5.509010000e-07 V_low
+ 5.510000000e-07 V_low
+ 5.510010000e-07 V_low
+ 5.511000000e-07 V_low
+ 5.511010000e-07 V_low
+ 5.512000000e-07 V_low
+ 5.512010000e-07 V_low
+ 5.513000000e-07 V_low
+ 5.513010000e-07 V_low
+ 5.514000000e-07 V_low
+ 5.514010000e-07 V_low
+ 5.515000000e-07 V_low
+ 5.515010000e-07 V_low
+ 5.516000000e-07 V_low
+ 5.516010000e-07 V_low
+ 5.517000000e-07 V_low
+ 5.517010000e-07 V_low
+ 5.518000000e-07 V_low
+ 5.518010000e-07 V_low
+ 5.519000000e-07 V_low
+ 5.519010000e-07 V_hig
+ 5.520000000e-07 V_hig
+ 5.520010000e-07 V_hig
+ 5.521000000e-07 V_hig
+ 5.521010000e-07 V_hig
+ 5.522000000e-07 V_hig
+ 5.522010000e-07 V_hig
+ 5.523000000e-07 V_hig
+ 5.523010000e-07 V_hig
+ 5.524000000e-07 V_hig
+ 5.524010000e-07 V_hig
+ 5.525000000e-07 V_hig
+ 5.525010000e-07 V_hig
+ 5.526000000e-07 V_hig
+ 5.526010000e-07 V_hig
+ 5.527000000e-07 V_hig
+ 5.527010000e-07 V_hig
+ 5.528000000e-07 V_hig
+ 5.528010000e-07 V_hig
+ 5.529000000e-07 V_hig
+ 5.529010000e-07 V_low
+ 5.530000000e-07 V_low
+ 5.530010000e-07 V_low
+ 5.531000000e-07 V_low
+ 5.531010000e-07 V_low
+ 5.532000000e-07 V_low
+ 5.532010000e-07 V_low
+ 5.533000000e-07 V_low
+ 5.533010000e-07 V_low
+ 5.534000000e-07 V_low
+ 5.534010000e-07 V_low
+ 5.535000000e-07 V_low
+ 5.535010000e-07 V_low
+ 5.536000000e-07 V_low
+ 5.536010000e-07 V_low
+ 5.537000000e-07 V_low
+ 5.537010000e-07 V_low
+ 5.538000000e-07 V_low
+ 5.538010000e-07 V_low
+ 5.539000000e-07 V_low
+ 5.539010000e-07 V_hig
+ 5.540000000e-07 V_hig
+ 5.540010000e-07 V_hig
+ 5.541000000e-07 V_hig
+ 5.541010000e-07 V_hig
+ 5.542000000e-07 V_hig
+ 5.542010000e-07 V_hig
+ 5.543000000e-07 V_hig
+ 5.543010000e-07 V_hig
+ 5.544000000e-07 V_hig
+ 5.544010000e-07 V_hig
+ 5.545000000e-07 V_hig
+ 5.545010000e-07 V_hig
+ 5.546000000e-07 V_hig
+ 5.546010000e-07 V_hig
+ 5.547000000e-07 V_hig
+ 5.547010000e-07 V_hig
+ 5.548000000e-07 V_hig
+ 5.548010000e-07 V_hig
+ 5.549000000e-07 V_hig
+ 5.549010000e-07 V_low
+ 5.550000000e-07 V_low
+ 5.550010000e-07 V_low
+ 5.551000000e-07 V_low
+ 5.551010000e-07 V_low
+ 5.552000000e-07 V_low
+ 5.552010000e-07 V_low
+ 5.553000000e-07 V_low
+ 5.553010000e-07 V_low
+ 5.554000000e-07 V_low
+ 5.554010000e-07 V_low
+ 5.555000000e-07 V_low
+ 5.555010000e-07 V_low
+ 5.556000000e-07 V_low
+ 5.556010000e-07 V_low
+ 5.557000000e-07 V_low
+ 5.557010000e-07 V_low
+ 5.558000000e-07 V_low
+ 5.558010000e-07 V_low
+ 5.559000000e-07 V_low
+ 5.559010000e-07 V_low
+ 5.560000000e-07 V_low
+ 5.560010000e-07 V_low
+ 5.561000000e-07 V_low
+ 5.561010000e-07 V_low
+ 5.562000000e-07 V_low
+ 5.562010000e-07 V_low
+ 5.563000000e-07 V_low
+ 5.563010000e-07 V_low
+ 5.564000000e-07 V_low
+ 5.564010000e-07 V_low
+ 5.565000000e-07 V_low
+ 5.565010000e-07 V_low
+ 5.566000000e-07 V_low
+ 5.566010000e-07 V_low
+ 5.567000000e-07 V_low
+ 5.567010000e-07 V_low
+ 5.568000000e-07 V_low
+ 5.568010000e-07 V_low
+ 5.569000000e-07 V_low
+ 5.569010000e-07 V_low
+ 5.570000000e-07 V_low
+ 5.570010000e-07 V_low
+ 5.571000000e-07 V_low
+ 5.571010000e-07 V_low
+ 5.572000000e-07 V_low
+ 5.572010000e-07 V_low
+ 5.573000000e-07 V_low
+ 5.573010000e-07 V_low
+ 5.574000000e-07 V_low
+ 5.574010000e-07 V_low
+ 5.575000000e-07 V_low
+ 5.575010000e-07 V_low
+ 5.576000000e-07 V_low
+ 5.576010000e-07 V_low
+ 5.577000000e-07 V_low
+ 5.577010000e-07 V_low
+ 5.578000000e-07 V_low
+ 5.578010000e-07 V_low
+ 5.579000000e-07 V_low
+ 5.579010000e-07 V_hig
+ 5.580000000e-07 V_hig
+ 5.580010000e-07 V_hig
+ 5.581000000e-07 V_hig
+ 5.581010000e-07 V_hig
+ 5.582000000e-07 V_hig
+ 5.582010000e-07 V_hig
+ 5.583000000e-07 V_hig
+ 5.583010000e-07 V_hig
+ 5.584000000e-07 V_hig
+ 5.584010000e-07 V_hig
+ 5.585000000e-07 V_hig
+ 5.585010000e-07 V_hig
+ 5.586000000e-07 V_hig
+ 5.586010000e-07 V_hig
+ 5.587000000e-07 V_hig
+ 5.587010000e-07 V_hig
+ 5.588000000e-07 V_hig
+ 5.588010000e-07 V_hig
+ 5.589000000e-07 V_hig
+ 5.589010000e-07 V_low
+ 5.590000000e-07 V_low
+ 5.590010000e-07 V_low
+ 5.591000000e-07 V_low
+ 5.591010000e-07 V_low
+ 5.592000000e-07 V_low
+ 5.592010000e-07 V_low
+ 5.593000000e-07 V_low
+ 5.593010000e-07 V_low
+ 5.594000000e-07 V_low
+ 5.594010000e-07 V_low
+ 5.595000000e-07 V_low
+ 5.595010000e-07 V_low
+ 5.596000000e-07 V_low
+ 5.596010000e-07 V_low
+ 5.597000000e-07 V_low
+ 5.597010000e-07 V_low
+ 5.598000000e-07 V_low
+ 5.598010000e-07 V_low
+ 5.599000000e-07 V_low
+ 5.599010000e-07 V_hig
+ 5.600000000e-07 V_hig
+ 5.600010000e-07 V_hig
+ 5.601000000e-07 V_hig
+ 5.601010000e-07 V_hig
+ 5.602000000e-07 V_hig
+ 5.602010000e-07 V_hig
+ 5.603000000e-07 V_hig
+ 5.603010000e-07 V_hig
+ 5.604000000e-07 V_hig
+ 5.604010000e-07 V_hig
+ 5.605000000e-07 V_hig
+ 5.605010000e-07 V_hig
+ 5.606000000e-07 V_hig
+ 5.606010000e-07 V_hig
+ 5.607000000e-07 V_hig
+ 5.607010000e-07 V_hig
+ 5.608000000e-07 V_hig
+ 5.608010000e-07 V_hig
+ 5.609000000e-07 V_hig
+ 5.609010000e-07 V_low
+ 5.610000000e-07 V_low
+ 5.610010000e-07 V_low
+ 5.611000000e-07 V_low
+ 5.611010000e-07 V_low
+ 5.612000000e-07 V_low
+ 5.612010000e-07 V_low
+ 5.613000000e-07 V_low
+ 5.613010000e-07 V_low
+ 5.614000000e-07 V_low
+ 5.614010000e-07 V_low
+ 5.615000000e-07 V_low
+ 5.615010000e-07 V_low
+ 5.616000000e-07 V_low
+ 5.616010000e-07 V_low
+ 5.617000000e-07 V_low
+ 5.617010000e-07 V_low
+ 5.618000000e-07 V_low
+ 5.618010000e-07 V_low
+ 5.619000000e-07 V_low
+ 5.619010000e-07 V_hig
+ 5.620000000e-07 V_hig
+ 5.620010000e-07 V_hig
+ 5.621000000e-07 V_hig
+ 5.621010000e-07 V_hig
+ 5.622000000e-07 V_hig
+ 5.622010000e-07 V_hig
+ 5.623000000e-07 V_hig
+ 5.623010000e-07 V_hig
+ 5.624000000e-07 V_hig
+ 5.624010000e-07 V_hig
+ 5.625000000e-07 V_hig
+ 5.625010000e-07 V_hig
+ 5.626000000e-07 V_hig
+ 5.626010000e-07 V_hig
+ 5.627000000e-07 V_hig
+ 5.627010000e-07 V_hig
+ 5.628000000e-07 V_hig
+ 5.628010000e-07 V_hig
+ 5.629000000e-07 V_hig
+ 5.629010000e-07 V_hig
+ 5.630000000e-07 V_hig
+ 5.630010000e-07 V_hig
+ 5.631000000e-07 V_hig
+ 5.631010000e-07 V_hig
+ 5.632000000e-07 V_hig
+ 5.632010000e-07 V_hig
+ 5.633000000e-07 V_hig
+ 5.633010000e-07 V_hig
+ 5.634000000e-07 V_hig
+ 5.634010000e-07 V_hig
+ 5.635000000e-07 V_hig
+ 5.635010000e-07 V_hig
+ 5.636000000e-07 V_hig
+ 5.636010000e-07 V_hig
+ 5.637000000e-07 V_hig
+ 5.637010000e-07 V_hig
+ 5.638000000e-07 V_hig
+ 5.638010000e-07 V_hig
+ 5.639000000e-07 V_hig
+ 5.639010000e-07 V_hig
+ 5.640000000e-07 V_hig
+ 5.640010000e-07 V_hig
+ 5.641000000e-07 V_hig
+ 5.641010000e-07 V_hig
+ 5.642000000e-07 V_hig
+ 5.642010000e-07 V_hig
+ 5.643000000e-07 V_hig
+ 5.643010000e-07 V_hig
+ 5.644000000e-07 V_hig
+ 5.644010000e-07 V_hig
+ 5.645000000e-07 V_hig
+ 5.645010000e-07 V_hig
+ 5.646000000e-07 V_hig
+ 5.646010000e-07 V_hig
+ 5.647000000e-07 V_hig
+ 5.647010000e-07 V_hig
+ 5.648000000e-07 V_hig
+ 5.648010000e-07 V_hig
+ 5.649000000e-07 V_hig
+ 5.649010000e-07 V_low
+ 5.650000000e-07 V_low
+ 5.650010000e-07 V_low
+ 5.651000000e-07 V_low
+ 5.651010000e-07 V_low
+ 5.652000000e-07 V_low
+ 5.652010000e-07 V_low
+ 5.653000000e-07 V_low
+ 5.653010000e-07 V_low
+ 5.654000000e-07 V_low
+ 5.654010000e-07 V_low
+ 5.655000000e-07 V_low
+ 5.655010000e-07 V_low
+ 5.656000000e-07 V_low
+ 5.656010000e-07 V_low
+ 5.657000000e-07 V_low
+ 5.657010000e-07 V_low
+ 5.658000000e-07 V_low
+ 5.658010000e-07 V_low
+ 5.659000000e-07 V_low
+ 5.659010000e-07 V_low
+ 5.660000000e-07 V_low
+ 5.660010000e-07 V_low
+ 5.661000000e-07 V_low
+ 5.661010000e-07 V_low
+ 5.662000000e-07 V_low
+ 5.662010000e-07 V_low
+ 5.663000000e-07 V_low
+ 5.663010000e-07 V_low
+ 5.664000000e-07 V_low
+ 5.664010000e-07 V_low
+ 5.665000000e-07 V_low
+ 5.665010000e-07 V_low
+ 5.666000000e-07 V_low
+ 5.666010000e-07 V_low
+ 5.667000000e-07 V_low
+ 5.667010000e-07 V_low
+ 5.668000000e-07 V_low
+ 5.668010000e-07 V_low
+ 5.669000000e-07 V_low
+ 5.669010000e-07 V_hig
+ 5.670000000e-07 V_hig
+ 5.670010000e-07 V_hig
+ 5.671000000e-07 V_hig
+ 5.671010000e-07 V_hig
+ 5.672000000e-07 V_hig
+ 5.672010000e-07 V_hig
+ 5.673000000e-07 V_hig
+ 5.673010000e-07 V_hig
+ 5.674000000e-07 V_hig
+ 5.674010000e-07 V_hig
+ 5.675000000e-07 V_hig
+ 5.675010000e-07 V_hig
+ 5.676000000e-07 V_hig
+ 5.676010000e-07 V_hig
+ 5.677000000e-07 V_hig
+ 5.677010000e-07 V_hig
+ 5.678000000e-07 V_hig
+ 5.678010000e-07 V_hig
+ 5.679000000e-07 V_hig
+ 5.679010000e-07 V_low
+ 5.680000000e-07 V_low
+ 5.680010000e-07 V_low
+ 5.681000000e-07 V_low
+ 5.681010000e-07 V_low
+ 5.682000000e-07 V_low
+ 5.682010000e-07 V_low
+ 5.683000000e-07 V_low
+ 5.683010000e-07 V_low
+ 5.684000000e-07 V_low
+ 5.684010000e-07 V_low
+ 5.685000000e-07 V_low
+ 5.685010000e-07 V_low
+ 5.686000000e-07 V_low
+ 5.686010000e-07 V_low
+ 5.687000000e-07 V_low
+ 5.687010000e-07 V_low
+ 5.688000000e-07 V_low
+ 5.688010000e-07 V_low
+ 5.689000000e-07 V_low
+ 5.689010000e-07 V_hig
+ 5.690000000e-07 V_hig
+ 5.690010000e-07 V_hig
+ 5.691000000e-07 V_hig
+ 5.691010000e-07 V_hig
+ 5.692000000e-07 V_hig
+ 5.692010000e-07 V_hig
+ 5.693000000e-07 V_hig
+ 5.693010000e-07 V_hig
+ 5.694000000e-07 V_hig
+ 5.694010000e-07 V_hig
+ 5.695000000e-07 V_hig
+ 5.695010000e-07 V_hig
+ 5.696000000e-07 V_hig
+ 5.696010000e-07 V_hig
+ 5.697000000e-07 V_hig
+ 5.697010000e-07 V_hig
+ 5.698000000e-07 V_hig
+ 5.698010000e-07 V_hig
+ 5.699000000e-07 V_hig
+ 5.699010000e-07 V_low
+ 5.700000000e-07 V_low
+ 5.700010000e-07 V_low
+ 5.701000000e-07 V_low
+ 5.701010000e-07 V_low
+ 5.702000000e-07 V_low
+ 5.702010000e-07 V_low
+ 5.703000000e-07 V_low
+ 5.703010000e-07 V_low
+ 5.704000000e-07 V_low
+ 5.704010000e-07 V_low
+ 5.705000000e-07 V_low
+ 5.705010000e-07 V_low
+ 5.706000000e-07 V_low
+ 5.706010000e-07 V_low
+ 5.707000000e-07 V_low
+ 5.707010000e-07 V_low
+ 5.708000000e-07 V_low
+ 5.708010000e-07 V_low
+ 5.709000000e-07 V_low
+ 5.709010000e-07 V_low
+ 5.710000000e-07 V_low
+ 5.710010000e-07 V_low
+ 5.711000000e-07 V_low
+ 5.711010000e-07 V_low
+ 5.712000000e-07 V_low
+ 5.712010000e-07 V_low
+ 5.713000000e-07 V_low
+ 5.713010000e-07 V_low
+ 5.714000000e-07 V_low
+ 5.714010000e-07 V_low
+ 5.715000000e-07 V_low
+ 5.715010000e-07 V_low
+ 5.716000000e-07 V_low
+ 5.716010000e-07 V_low
+ 5.717000000e-07 V_low
+ 5.717010000e-07 V_low
+ 5.718000000e-07 V_low
+ 5.718010000e-07 V_low
+ 5.719000000e-07 V_low
+ 5.719010000e-07 V_low
+ 5.720000000e-07 V_low
+ 5.720010000e-07 V_low
+ 5.721000000e-07 V_low
+ 5.721010000e-07 V_low
+ 5.722000000e-07 V_low
+ 5.722010000e-07 V_low
+ 5.723000000e-07 V_low
+ 5.723010000e-07 V_low
+ 5.724000000e-07 V_low
+ 5.724010000e-07 V_low
+ 5.725000000e-07 V_low
+ 5.725010000e-07 V_low
+ 5.726000000e-07 V_low
+ 5.726010000e-07 V_low
+ 5.727000000e-07 V_low
+ 5.727010000e-07 V_low
+ 5.728000000e-07 V_low
+ 5.728010000e-07 V_low
+ 5.729000000e-07 V_low
+ 5.729010000e-07 V_hig
+ 5.730000000e-07 V_hig
+ 5.730010000e-07 V_hig
+ 5.731000000e-07 V_hig
+ 5.731010000e-07 V_hig
+ 5.732000000e-07 V_hig
+ 5.732010000e-07 V_hig
+ 5.733000000e-07 V_hig
+ 5.733010000e-07 V_hig
+ 5.734000000e-07 V_hig
+ 5.734010000e-07 V_hig
+ 5.735000000e-07 V_hig
+ 5.735010000e-07 V_hig
+ 5.736000000e-07 V_hig
+ 5.736010000e-07 V_hig
+ 5.737000000e-07 V_hig
+ 5.737010000e-07 V_hig
+ 5.738000000e-07 V_hig
+ 5.738010000e-07 V_hig
+ 5.739000000e-07 V_hig
+ 5.739010000e-07 V_hig
+ 5.740000000e-07 V_hig
+ 5.740010000e-07 V_hig
+ 5.741000000e-07 V_hig
+ 5.741010000e-07 V_hig
+ 5.742000000e-07 V_hig
+ 5.742010000e-07 V_hig
+ 5.743000000e-07 V_hig
+ 5.743010000e-07 V_hig
+ 5.744000000e-07 V_hig
+ 5.744010000e-07 V_hig
+ 5.745000000e-07 V_hig
+ 5.745010000e-07 V_hig
+ 5.746000000e-07 V_hig
+ 5.746010000e-07 V_hig
+ 5.747000000e-07 V_hig
+ 5.747010000e-07 V_hig
+ 5.748000000e-07 V_hig
+ 5.748010000e-07 V_hig
+ 5.749000000e-07 V_hig
+ 5.749010000e-07 V_hig
+ 5.750000000e-07 V_hig
+ 5.750010000e-07 V_hig
+ 5.751000000e-07 V_hig
+ 5.751010000e-07 V_hig
+ 5.752000000e-07 V_hig
+ 5.752010000e-07 V_hig
+ 5.753000000e-07 V_hig
+ 5.753010000e-07 V_hig
+ 5.754000000e-07 V_hig
+ 5.754010000e-07 V_hig
+ 5.755000000e-07 V_hig
+ 5.755010000e-07 V_hig
+ 5.756000000e-07 V_hig
+ 5.756010000e-07 V_hig
+ 5.757000000e-07 V_hig
+ 5.757010000e-07 V_hig
+ 5.758000000e-07 V_hig
+ 5.758010000e-07 V_hig
+ 5.759000000e-07 V_hig
+ 5.759010000e-07 V_low
+ 5.760000000e-07 V_low
+ 5.760010000e-07 V_low
+ 5.761000000e-07 V_low
+ 5.761010000e-07 V_low
+ 5.762000000e-07 V_low
+ 5.762010000e-07 V_low
+ 5.763000000e-07 V_low
+ 5.763010000e-07 V_low
+ 5.764000000e-07 V_low
+ 5.764010000e-07 V_low
+ 5.765000000e-07 V_low
+ 5.765010000e-07 V_low
+ 5.766000000e-07 V_low
+ 5.766010000e-07 V_low
+ 5.767000000e-07 V_low
+ 5.767010000e-07 V_low
+ 5.768000000e-07 V_low
+ 5.768010000e-07 V_low
+ 5.769000000e-07 V_low
+ 5.769010000e-07 V_low
+ 5.770000000e-07 V_low
+ 5.770010000e-07 V_low
+ 5.771000000e-07 V_low
+ 5.771010000e-07 V_low
+ 5.772000000e-07 V_low
+ 5.772010000e-07 V_low
+ 5.773000000e-07 V_low
+ 5.773010000e-07 V_low
+ 5.774000000e-07 V_low
+ 5.774010000e-07 V_low
+ 5.775000000e-07 V_low
+ 5.775010000e-07 V_low
+ 5.776000000e-07 V_low
+ 5.776010000e-07 V_low
+ 5.777000000e-07 V_low
+ 5.777010000e-07 V_low
+ 5.778000000e-07 V_low
+ 5.778010000e-07 V_low
+ 5.779000000e-07 V_low
+ 5.779010000e-07 V_low
+ 5.780000000e-07 V_low
+ 5.780010000e-07 V_low
+ 5.781000000e-07 V_low
+ 5.781010000e-07 V_low
+ 5.782000000e-07 V_low
+ 5.782010000e-07 V_low
+ 5.783000000e-07 V_low
+ 5.783010000e-07 V_low
+ 5.784000000e-07 V_low
+ 5.784010000e-07 V_low
+ 5.785000000e-07 V_low
+ 5.785010000e-07 V_low
+ 5.786000000e-07 V_low
+ 5.786010000e-07 V_low
+ 5.787000000e-07 V_low
+ 5.787010000e-07 V_low
+ 5.788000000e-07 V_low
+ 5.788010000e-07 V_low
+ 5.789000000e-07 V_low
+ 5.789010000e-07 V_hig
+ 5.790000000e-07 V_hig
+ 5.790010000e-07 V_hig
+ 5.791000000e-07 V_hig
+ 5.791010000e-07 V_hig
+ 5.792000000e-07 V_hig
+ 5.792010000e-07 V_hig
+ 5.793000000e-07 V_hig
+ 5.793010000e-07 V_hig
+ 5.794000000e-07 V_hig
+ 5.794010000e-07 V_hig
+ 5.795000000e-07 V_hig
+ 5.795010000e-07 V_hig
+ 5.796000000e-07 V_hig
+ 5.796010000e-07 V_hig
+ 5.797000000e-07 V_hig
+ 5.797010000e-07 V_hig
+ 5.798000000e-07 V_hig
+ 5.798010000e-07 V_hig
+ 5.799000000e-07 V_hig
+ 5.799010000e-07 V_low
+ 5.800000000e-07 V_low
+ 5.800010000e-07 V_low
+ 5.801000000e-07 V_low
+ 5.801010000e-07 V_low
+ 5.802000000e-07 V_low
+ 5.802010000e-07 V_low
+ 5.803000000e-07 V_low
+ 5.803010000e-07 V_low
+ 5.804000000e-07 V_low
+ 5.804010000e-07 V_low
+ 5.805000000e-07 V_low
+ 5.805010000e-07 V_low
+ 5.806000000e-07 V_low
+ 5.806010000e-07 V_low
+ 5.807000000e-07 V_low
+ 5.807010000e-07 V_low
+ 5.808000000e-07 V_low
+ 5.808010000e-07 V_low
+ 5.809000000e-07 V_low
+ 5.809010000e-07 V_hig
+ 5.810000000e-07 V_hig
+ 5.810010000e-07 V_hig
+ 5.811000000e-07 V_hig
+ 5.811010000e-07 V_hig
+ 5.812000000e-07 V_hig
+ 5.812010000e-07 V_hig
+ 5.813000000e-07 V_hig
+ 5.813010000e-07 V_hig
+ 5.814000000e-07 V_hig
+ 5.814010000e-07 V_hig
+ 5.815000000e-07 V_hig
+ 5.815010000e-07 V_hig
+ 5.816000000e-07 V_hig
+ 5.816010000e-07 V_hig
+ 5.817000000e-07 V_hig
+ 5.817010000e-07 V_hig
+ 5.818000000e-07 V_hig
+ 5.818010000e-07 V_hig
+ 5.819000000e-07 V_hig
+ 5.819010000e-07 V_hig
+ 5.820000000e-07 V_hig
+ 5.820010000e-07 V_hig
+ 5.821000000e-07 V_hig
+ 5.821010000e-07 V_hig
+ 5.822000000e-07 V_hig
+ 5.822010000e-07 V_hig
+ 5.823000000e-07 V_hig
+ 5.823010000e-07 V_hig
+ 5.824000000e-07 V_hig
+ 5.824010000e-07 V_hig
+ 5.825000000e-07 V_hig
+ 5.825010000e-07 V_hig
+ 5.826000000e-07 V_hig
+ 5.826010000e-07 V_hig
+ 5.827000000e-07 V_hig
+ 5.827010000e-07 V_hig
+ 5.828000000e-07 V_hig
+ 5.828010000e-07 V_hig
+ 5.829000000e-07 V_hig
+ 5.829010000e-07 V_low
+ 5.830000000e-07 V_low
+ 5.830010000e-07 V_low
+ 5.831000000e-07 V_low
+ 5.831010000e-07 V_low
+ 5.832000000e-07 V_low
+ 5.832010000e-07 V_low
+ 5.833000000e-07 V_low
+ 5.833010000e-07 V_low
+ 5.834000000e-07 V_low
+ 5.834010000e-07 V_low
+ 5.835000000e-07 V_low
+ 5.835010000e-07 V_low
+ 5.836000000e-07 V_low
+ 5.836010000e-07 V_low
+ 5.837000000e-07 V_low
+ 5.837010000e-07 V_low
+ 5.838000000e-07 V_low
+ 5.838010000e-07 V_low
+ 5.839000000e-07 V_low
+ 5.839010000e-07 V_low
+ 5.840000000e-07 V_low
+ 5.840010000e-07 V_low
+ 5.841000000e-07 V_low
+ 5.841010000e-07 V_low
+ 5.842000000e-07 V_low
+ 5.842010000e-07 V_low
+ 5.843000000e-07 V_low
+ 5.843010000e-07 V_low
+ 5.844000000e-07 V_low
+ 5.844010000e-07 V_low
+ 5.845000000e-07 V_low
+ 5.845010000e-07 V_low
+ 5.846000000e-07 V_low
+ 5.846010000e-07 V_low
+ 5.847000000e-07 V_low
+ 5.847010000e-07 V_low
+ 5.848000000e-07 V_low
+ 5.848010000e-07 V_low
+ 5.849000000e-07 V_low
+ 5.849010000e-07 V_hig
+ 5.850000000e-07 V_hig
+ 5.850010000e-07 V_hig
+ 5.851000000e-07 V_hig
+ 5.851010000e-07 V_hig
+ 5.852000000e-07 V_hig
+ 5.852010000e-07 V_hig
+ 5.853000000e-07 V_hig
+ 5.853010000e-07 V_hig
+ 5.854000000e-07 V_hig
+ 5.854010000e-07 V_hig
+ 5.855000000e-07 V_hig
+ 5.855010000e-07 V_hig
+ 5.856000000e-07 V_hig
+ 5.856010000e-07 V_hig
+ 5.857000000e-07 V_hig
+ 5.857010000e-07 V_hig
+ 5.858000000e-07 V_hig
+ 5.858010000e-07 V_hig
+ 5.859000000e-07 V_hig
+ 5.859010000e-07 V_hig
+ 5.860000000e-07 V_hig
+ 5.860010000e-07 V_hig
+ 5.861000000e-07 V_hig
+ 5.861010000e-07 V_hig
+ 5.862000000e-07 V_hig
+ 5.862010000e-07 V_hig
+ 5.863000000e-07 V_hig
+ 5.863010000e-07 V_hig
+ 5.864000000e-07 V_hig
+ 5.864010000e-07 V_hig
+ 5.865000000e-07 V_hig
+ 5.865010000e-07 V_hig
+ 5.866000000e-07 V_hig
+ 5.866010000e-07 V_hig
+ 5.867000000e-07 V_hig
+ 5.867010000e-07 V_hig
+ 5.868000000e-07 V_hig
+ 5.868010000e-07 V_hig
+ 5.869000000e-07 V_hig
+ 5.869010000e-07 V_low
+ 5.870000000e-07 V_low
+ 5.870010000e-07 V_low
+ 5.871000000e-07 V_low
+ 5.871010000e-07 V_low
+ 5.872000000e-07 V_low
+ 5.872010000e-07 V_low
+ 5.873000000e-07 V_low
+ 5.873010000e-07 V_low
+ 5.874000000e-07 V_low
+ 5.874010000e-07 V_low
+ 5.875000000e-07 V_low
+ 5.875010000e-07 V_low
+ 5.876000000e-07 V_low
+ 5.876010000e-07 V_low
+ 5.877000000e-07 V_low
+ 5.877010000e-07 V_low
+ 5.878000000e-07 V_low
+ 5.878010000e-07 V_low
+ 5.879000000e-07 V_low
+ 5.879010000e-07 V_hig
+ 5.880000000e-07 V_hig
+ 5.880010000e-07 V_hig
+ 5.881000000e-07 V_hig
+ 5.881010000e-07 V_hig
+ 5.882000000e-07 V_hig
+ 5.882010000e-07 V_hig
+ 5.883000000e-07 V_hig
+ 5.883010000e-07 V_hig
+ 5.884000000e-07 V_hig
+ 5.884010000e-07 V_hig
+ 5.885000000e-07 V_hig
+ 5.885010000e-07 V_hig
+ 5.886000000e-07 V_hig
+ 5.886010000e-07 V_hig
+ 5.887000000e-07 V_hig
+ 5.887010000e-07 V_hig
+ 5.888000000e-07 V_hig
+ 5.888010000e-07 V_hig
+ 5.889000000e-07 V_hig
+ 5.889010000e-07 V_hig
+ 5.890000000e-07 V_hig
+ 5.890010000e-07 V_hig
+ 5.891000000e-07 V_hig
+ 5.891010000e-07 V_hig
+ 5.892000000e-07 V_hig
+ 5.892010000e-07 V_hig
+ 5.893000000e-07 V_hig
+ 5.893010000e-07 V_hig
+ 5.894000000e-07 V_hig
+ 5.894010000e-07 V_hig
+ 5.895000000e-07 V_hig
+ 5.895010000e-07 V_hig
+ 5.896000000e-07 V_hig
+ 5.896010000e-07 V_hig
+ 5.897000000e-07 V_hig
+ 5.897010000e-07 V_hig
+ 5.898000000e-07 V_hig
+ 5.898010000e-07 V_hig
+ 5.899000000e-07 V_hig
+ 5.899010000e-07 V_hig
+ 5.900000000e-07 V_hig
+ 5.900010000e-07 V_hig
+ 5.901000000e-07 V_hig
+ 5.901010000e-07 V_hig
+ 5.902000000e-07 V_hig
+ 5.902010000e-07 V_hig
+ 5.903000000e-07 V_hig
+ 5.903010000e-07 V_hig
+ 5.904000000e-07 V_hig
+ 5.904010000e-07 V_hig
+ 5.905000000e-07 V_hig
+ 5.905010000e-07 V_hig
+ 5.906000000e-07 V_hig
+ 5.906010000e-07 V_hig
+ 5.907000000e-07 V_hig
+ 5.907010000e-07 V_hig
+ 5.908000000e-07 V_hig
+ 5.908010000e-07 V_hig
+ 5.909000000e-07 V_hig
+ 5.909010000e-07 V_low
+ 5.910000000e-07 V_low
+ 5.910010000e-07 V_low
+ 5.911000000e-07 V_low
+ 5.911010000e-07 V_low
+ 5.912000000e-07 V_low
+ 5.912010000e-07 V_low
+ 5.913000000e-07 V_low
+ 5.913010000e-07 V_low
+ 5.914000000e-07 V_low
+ 5.914010000e-07 V_low
+ 5.915000000e-07 V_low
+ 5.915010000e-07 V_low
+ 5.916000000e-07 V_low
+ 5.916010000e-07 V_low
+ 5.917000000e-07 V_low
+ 5.917010000e-07 V_low
+ 5.918000000e-07 V_low
+ 5.918010000e-07 V_low
+ 5.919000000e-07 V_low
+ 5.919010000e-07 V_hig
+ 5.920000000e-07 V_hig
+ 5.920010000e-07 V_hig
+ 5.921000000e-07 V_hig
+ 5.921010000e-07 V_hig
+ 5.922000000e-07 V_hig
+ 5.922010000e-07 V_hig
+ 5.923000000e-07 V_hig
+ 5.923010000e-07 V_hig
+ 5.924000000e-07 V_hig
+ 5.924010000e-07 V_hig
+ 5.925000000e-07 V_hig
+ 5.925010000e-07 V_hig
+ 5.926000000e-07 V_hig
+ 5.926010000e-07 V_hig
+ 5.927000000e-07 V_hig
+ 5.927010000e-07 V_hig
+ 5.928000000e-07 V_hig
+ 5.928010000e-07 V_hig
+ 5.929000000e-07 V_hig
+ 5.929010000e-07 V_low
+ 5.930000000e-07 V_low
+ 5.930010000e-07 V_low
+ 5.931000000e-07 V_low
+ 5.931010000e-07 V_low
+ 5.932000000e-07 V_low
+ 5.932010000e-07 V_low
+ 5.933000000e-07 V_low
+ 5.933010000e-07 V_low
+ 5.934000000e-07 V_low
+ 5.934010000e-07 V_low
+ 5.935000000e-07 V_low
+ 5.935010000e-07 V_low
+ 5.936000000e-07 V_low
+ 5.936010000e-07 V_low
+ 5.937000000e-07 V_low
+ 5.937010000e-07 V_low
+ 5.938000000e-07 V_low
+ 5.938010000e-07 V_low
+ 5.939000000e-07 V_low
+ 5.939010000e-07 V_hig
+ 5.940000000e-07 V_hig
+ 5.940010000e-07 V_hig
+ 5.941000000e-07 V_hig
+ 5.941010000e-07 V_hig
+ 5.942000000e-07 V_hig
+ 5.942010000e-07 V_hig
+ 5.943000000e-07 V_hig
+ 5.943010000e-07 V_hig
+ 5.944000000e-07 V_hig
+ 5.944010000e-07 V_hig
+ 5.945000000e-07 V_hig
+ 5.945010000e-07 V_hig
+ 5.946000000e-07 V_hig
+ 5.946010000e-07 V_hig
+ 5.947000000e-07 V_hig
+ 5.947010000e-07 V_hig
+ 5.948000000e-07 V_hig
+ 5.948010000e-07 V_hig
+ 5.949000000e-07 V_hig
+ 5.949010000e-07 V_hig
+ 5.950000000e-07 V_hig
+ 5.950010000e-07 V_hig
+ 5.951000000e-07 V_hig
+ 5.951010000e-07 V_hig
+ 5.952000000e-07 V_hig
+ 5.952010000e-07 V_hig
+ 5.953000000e-07 V_hig
+ 5.953010000e-07 V_hig
+ 5.954000000e-07 V_hig
+ 5.954010000e-07 V_hig
+ 5.955000000e-07 V_hig
+ 5.955010000e-07 V_hig
+ 5.956000000e-07 V_hig
+ 5.956010000e-07 V_hig
+ 5.957000000e-07 V_hig
+ 5.957010000e-07 V_hig
+ 5.958000000e-07 V_hig
+ 5.958010000e-07 V_hig
+ 5.959000000e-07 V_hig
+ 5.959010000e-07 V_hig
+ 5.960000000e-07 V_hig
+ 5.960010000e-07 V_hig
+ 5.961000000e-07 V_hig
+ 5.961010000e-07 V_hig
+ 5.962000000e-07 V_hig
+ 5.962010000e-07 V_hig
+ 5.963000000e-07 V_hig
+ 5.963010000e-07 V_hig
+ 5.964000000e-07 V_hig
+ 5.964010000e-07 V_hig
+ 5.965000000e-07 V_hig
+ 5.965010000e-07 V_hig
+ 5.966000000e-07 V_hig
+ 5.966010000e-07 V_hig
+ 5.967000000e-07 V_hig
+ 5.967010000e-07 V_hig
+ 5.968000000e-07 V_hig
+ 5.968010000e-07 V_hig
+ 5.969000000e-07 V_hig
+ 5.969010000e-07 V_low
+ 5.970000000e-07 V_low
+ 5.970010000e-07 V_low
+ 5.971000000e-07 V_low
+ 5.971010000e-07 V_low
+ 5.972000000e-07 V_low
+ 5.972010000e-07 V_low
+ 5.973000000e-07 V_low
+ 5.973010000e-07 V_low
+ 5.974000000e-07 V_low
+ 5.974010000e-07 V_low
+ 5.975000000e-07 V_low
+ 5.975010000e-07 V_low
+ 5.976000000e-07 V_low
+ 5.976010000e-07 V_low
+ 5.977000000e-07 V_low
+ 5.977010000e-07 V_low
+ 5.978000000e-07 V_low
+ 5.978010000e-07 V_low
+ 5.979000000e-07 V_low
+ 5.979010000e-07 V_low
+ 5.980000000e-07 V_low
+ 5.980010000e-07 V_low
+ 5.981000000e-07 V_low
+ 5.981010000e-07 V_low
+ 5.982000000e-07 V_low
+ 5.982010000e-07 V_low
+ 5.983000000e-07 V_low
+ 5.983010000e-07 V_low
+ 5.984000000e-07 V_low
+ 5.984010000e-07 V_low
+ 5.985000000e-07 V_low
+ 5.985010000e-07 V_low
+ 5.986000000e-07 V_low
+ 5.986010000e-07 V_low
+ 5.987000000e-07 V_low
+ 5.987010000e-07 V_low
+ 5.988000000e-07 V_low
+ 5.988010000e-07 V_low
+ 5.989000000e-07 V_low
+ 5.989010000e-07 V_hig
+ 5.990000000e-07 V_hig
+ 5.990010000e-07 V_hig
+ 5.991000000e-07 V_hig
+ 5.991010000e-07 V_hig
+ 5.992000000e-07 V_hig
+ 5.992010000e-07 V_hig
+ 5.993000000e-07 V_hig
+ 5.993010000e-07 V_hig
+ 5.994000000e-07 V_hig
+ 5.994010000e-07 V_hig
+ 5.995000000e-07 V_hig
+ 5.995010000e-07 V_hig
+ 5.996000000e-07 V_hig
+ 5.996010000e-07 V_hig
+ 5.997000000e-07 V_hig
+ 5.997010000e-07 V_hig
+ 5.998000000e-07 V_hig
+ 5.998010000e-07 V_hig
+ 5.999000000e-07 V_hig
+ 5.999010000e-07 V_low
+ 6.000000000e-07 V_low
+ 6.000010000e-07 V_low
+ 6.001000000e-07 V_low
+ 6.001010000e-07 V_low
+ 6.002000000e-07 V_low
+ 6.002010000e-07 V_low
+ 6.003000000e-07 V_low
+ 6.003010000e-07 V_low
+ 6.004000000e-07 V_low
+ 6.004010000e-07 V_low
+ 6.005000000e-07 V_low
+ 6.005010000e-07 V_low
+ 6.006000000e-07 V_low
+ 6.006010000e-07 V_low
+ 6.007000000e-07 V_low
+ 6.007010000e-07 V_low
+ 6.008000000e-07 V_low
+ 6.008010000e-07 V_low
+ 6.009000000e-07 V_low
+ 6.009010000e-07 V_low
+ 6.010000000e-07 V_low
+ 6.010010000e-07 V_low
+ 6.011000000e-07 V_low
+ 6.011010000e-07 V_low
+ 6.012000000e-07 V_low
+ 6.012010000e-07 V_low
+ 6.013000000e-07 V_low
+ 6.013010000e-07 V_low
+ 6.014000000e-07 V_low
+ 6.014010000e-07 V_low
+ 6.015000000e-07 V_low
+ 6.015010000e-07 V_low
+ 6.016000000e-07 V_low
+ 6.016010000e-07 V_low
+ 6.017000000e-07 V_low
+ 6.017010000e-07 V_low
+ 6.018000000e-07 V_low
+ 6.018010000e-07 V_low
+ 6.019000000e-07 V_low
+ 6.019010000e-07 V_low
+ 6.020000000e-07 V_low
+ 6.020010000e-07 V_low
+ 6.021000000e-07 V_low
+ 6.021010000e-07 V_low
+ 6.022000000e-07 V_low
+ 6.022010000e-07 V_low
+ 6.023000000e-07 V_low
+ 6.023010000e-07 V_low
+ 6.024000000e-07 V_low
+ 6.024010000e-07 V_low
+ 6.025000000e-07 V_low
+ 6.025010000e-07 V_low
+ 6.026000000e-07 V_low
+ 6.026010000e-07 V_low
+ 6.027000000e-07 V_low
+ 6.027010000e-07 V_low
+ 6.028000000e-07 V_low
+ 6.028010000e-07 V_low
+ 6.029000000e-07 V_low
+ 6.029010000e-07 V_hig
+ 6.030000000e-07 V_hig
+ 6.030010000e-07 V_hig
+ 6.031000000e-07 V_hig
+ 6.031010000e-07 V_hig
+ 6.032000000e-07 V_hig
+ 6.032010000e-07 V_hig
+ 6.033000000e-07 V_hig
+ 6.033010000e-07 V_hig
+ 6.034000000e-07 V_hig
+ 6.034010000e-07 V_hig
+ 6.035000000e-07 V_hig
+ 6.035010000e-07 V_hig
+ 6.036000000e-07 V_hig
+ 6.036010000e-07 V_hig
+ 6.037000000e-07 V_hig
+ 6.037010000e-07 V_hig
+ 6.038000000e-07 V_hig
+ 6.038010000e-07 V_hig
+ 6.039000000e-07 V_hig
+ 6.039010000e-07 V_low
+ 6.040000000e-07 V_low
+ 6.040010000e-07 V_low
+ 6.041000000e-07 V_low
+ 6.041010000e-07 V_low
+ 6.042000000e-07 V_low
+ 6.042010000e-07 V_low
+ 6.043000000e-07 V_low
+ 6.043010000e-07 V_low
+ 6.044000000e-07 V_low
+ 6.044010000e-07 V_low
+ 6.045000000e-07 V_low
+ 6.045010000e-07 V_low
+ 6.046000000e-07 V_low
+ 6.046010000e-07 V_low
+ 6.047000000e-07 V_low
+ 6.047010000e-07 V_low
+ 6.048000000e-07 V_low
+ 6.048010000e-07 V_low
+ 6.049000000e-07 V_low
+ 6.049010000e-07 V_low
+ 6.050000000e-07 V_low
+ 6.050010000e-07 V_low
+ 6.051000000e-07 V_low
+ 6.051010000e-07 V_low
+ 6.052000000e-07 V_low
+ 6.052010000e-07 V_low
+ 6.053000000e-07 V_low
+ 6.053010000e-07 V_low
+ 6.054000000e-07 V_low
+ 6.054010000e-07 V_low
+ 6.055000000e-07 V_low
+ 6.055010000e-07 V_low
+ 6.056000000e-07 V_low
+ 6.056010000e-07 V_low
+ 6.057000000e-07 V_low
+ 6.057010000e-07 V_low
+ 6.058000000e-07 V_low
+ 6.058010000e-07 V_low
+ 6.059000000e-07 V_low
+ 6.059010000e-07 V_hig
+ 6.060000000e-07 V_hig
+ 6.060010000e-07 V_hig
+ 6.061000000e-07 V_hig
+ 6.061010000e-07 V_hig
+ 6.062000000e-07 V_hig
+ 6.062010000e-07 V_hig
+ 6.063000000e-07 V_hig
+ 6.063010000e-07 V_hig
+ 6.064000000e-07 V_hig
+ 6.064010000e-07 V_hig
+ 6.065000000e-07 V_hig
+ 6.065010000e-07 V_hig
+ 6.066000000e-07 V_hig
+ 6.066010000e-07 V_hig
+ 6.067000000e-07 V_hig
+ 6.067010000e-07 V_hig
+ 6.068000000e-07 V_hig
+ 6.068010000e-07 V_hig
+ 6.069000000e-07 V_hig
+ 6.069010000e-07 V_hig
+ 6.070000000e-07 V_hig
+ 6.070010000e-07 V_hig
+ 6.071000000e-07 V_hig
+ 6.071010000e-07 V_hig
+ 6.072000000e-07 V_hig
+ 6.072010000e-07 V_hig
+ 6.073000000e-07 V_hig
+ 6.073010000e-07 V_hig
+ 6.074000000e-07 V_hig
+ 6.074010000e-07 V_hig
+ 6.075000000e-07 V_hig
+ 6.075010000e-07 V_hig
+ 6.076000000e-07 V_hig
+ 6.076010000e-07 V_hig
+ 6.077000000e-07 V_hig
+ 6.077010000e-07 V_hig
+ 6.078000000e-07 V_hig
+ 6.078010000e-07 V_hig
+ 6.079000000e-07 V_hig
+ 6.079010000e-07 V_hig
+ 6.080000000e-07 V_hig
+ 6.080010000e-07 V_hig
+ 6.081000000e-07 V_hig
+ 6.081010000e-07 V_hig
+ 6.082000000e-07 V_hig
+ 6.082010000e-07 V_hig
+ 6.083000000e-07 V_hig
+ 6.083010000e-07 V_hig
+ 6.084000000e-07 V_hig
+ 6.084010000e-07 V_hig
+ 6.085000000e-07 V_hig
+ 6.085010000e-07 V_hig
+ 6.086000000e-07 V_hig
+ 6.086010000e-07 V_hig
+ 6.087000000e-07 V_hig
+ 6.087010000e-07 V_hig
+ 6.088000000e-07 V_hig
+ 6.088010000e-07 V_hig
+ 6.089000000e-07 V_hig
+ 6.089010000e-07 V_hig
+ 6.090000000e-07 V_hig
+ 6.090010000e-07 V_hig
+ 6.091000000e-07 V_hig
+ 6.091010000e-07 V_hig
+ 6.092000000e-07 V_hig
+ 6.092010000e-07 V_hig
+ 6.093000000e-07 V_hig
+ 6.093010000e-07 V_hig
+ 6.094000000e-07 V_hig
+ 6.094010000e-07 V_hig
+ 6.095000000e-07 V_hig
+ 6.095010000e-07 V_hig
+ 6.096000000e-07 V_hig
+ 6.096010000e-07 V_hig
+ 6.097000000e-07 V_hig
+ 6.097010000e-07 V_hig
+ 6.098000000e-07 V_hig
+ 6.098010000e-07 V_hig
+ 6.099000000e-07 V_hig
+ 6.099010000e-07 V_low
+ 6.100000000e-07 V_low
+ 6.100010000e-07 V_low
+ 6.101000000e-07 V_low
+ 6.101010000e-07 V_low
+ 6.102000000e-07 V_low
+ 6.102010000e-07 V_low
+ 6.103000000e-07 V_low
+ 6.103010000e-07 V_low
+ 6.104000000e-07 V_low
+ 6.104010000e-07 V_low
+ 6.105000000e-07 V_low
+ 6.105010000e-07 V_low
+ 6.106000000e-07 V_low
+ 6.106010000e-07 V_low
+ 6.107000000e-07 V_low
+ 6.107010000e-07 V_low
+ 6.108000000e-07 V_low
+ 6.108010000e-07 V_low
+ 6.109000000e-07 V_low
+ 6.109010000e-07 V_low
+ 6.110000000e-07 V_low
+ 6.110010000e-07 V_low
+ 6.111000000e-07 V_low
+ 6.111010000e-07 V_low
+ 6.112000000e-07 V_low
+ 6.112010000e-07 V_low
+ 6.113000000e-07 V_low
+ 6.113010000e-07 V_low
+ 6.114000000e-07 V_low
+ 6.114010000e-07 V_low
+ 6.115000000e-07 V_low
+ 6.115010000e-07 V_low
+ 6.116000000e-07 V_low
+ 6.116010000e-07 V_low
+ 6.117000000e-07 V_low
+ 6.117010000e-07 V_low
+ 6.118000000e-07 V_low
+ 6.118010000e-07 V_low
+ 6.119000000e-07 V_low
+ 6.119010000e-07 V_low
+ 6.120000000e-07 V_low
+ 6.120010000e-07 V_low
+ 6.121000000e-07 V_low
+ 6.121010000e-07 V_low
+ 6.122000000e-07 V_low
+ 6.122010000e-07 V_low
+ 6.123000000e-07 V_low
+ 6.123010000e-07 V_low
+ 6.124000000e-07 V_low
+ 6.124010000e-07 V_low
+ 6.125000000e-07 V_low
+ 6.125010000e-07 V_low
+ 6.126000000e-07 V_low
+ 6.126010000e-07 V_low
+ 6.127000000e-07 V_low
+ 6.127010000e-07 V_low
+ 6.128000000e-07 V_low
+ 6.128010000e-07 V_low
+ 6.129000000e-07 V_low
+ 6.129010000e-07 V_low
+ 6.130000000e-07 V_low
+ 6.130010000e-07 V_low
+ 6.131000000e-07 V_low
+ 6.131010000e-07 V_low
+ 6.132000000e-07 V_low
+ 6.132010000e-07 V_low
+ 6.133000000e-07 V_low
+ 6.133010000e-07 V_low
+ 6.134000000e-07 V_low
+ 6.134010000e-07 V_low
+ 6.135000000e-07 V_low
+ 6.135010000e-07 V_low
+ 6.136000000e-07 V_low
+ 6.136010000e-07 V_low
+ 6.137000000e-07 V_low
+ 6.137010000e-07 V_low
+ 6.138000000e-07 V_low
+ 6.138010000e-07 V_low
+ 6.139000000e-07 V_low
+ 6.139010000e-07 V_low
+ 6.140000000e-07 V_low
+ 6.140010000e-07 V_low
+ 6.141000000e-07 V_low
+ 6.141010000e-07 V_low
+ 6.142000000e-07 V_low
+ 6.142010000e-07 V_low
+ 6.143000000e-07 V_low
+ 6.143010000e-07 V_low
+ 6.144000000e-07 V_low
+ 6.144010000e-07 V_low
+ 6.145000000e-07 V_low
+ 6.145010000e-07 V_low
+ 6.146000000e-07 V_low
+ 6.146010000e-07 V_low
+ 6.147000000e-07 V_low
+ 6.147010000e-07 V_low
+ 6.148000000e-07 V_low
+ 6.148010000e-07 V_low
+ 6.149000000e-07 V_low
+ 6.149010000e-07 V_low
+ 6.150000000e-07 V_low
+ 6.150010000e-07 V_low
+ 6.151000000e-07 V_low
+ 6.151010000e-07 V_low
+ 6.152000000e-07 V_low
+ 6.152010000e-07 V_low
+ 6.153000000e-07 V_low
+ 6.153010000e-07 V_low
+ 6.154000000e-07 V_low
+ 6.154010000e-07 V_low
+ 6.155000000e-07 V_low
+ 6.155010000e-07 V_low
+ 6.156000000e-07 V_low
+ 6.156010000e-07 V_low
+ 6.157000000e-07 V_low
+ 6.157010000e-07 V_low
+ 6.158000000e-07 V_low
+ 6.158010000e-07 V_low
+ 6.159000000e-07 V_low
+ 6.159010000e-07 V_low
+ 6.160000000e-07 V_low
+ 6.160010000e-07 V_low
+ 6.161000000e-07 V_low
+ 6.161010000e-07 V_low
+ 6.162000000e-07 V_low
+ 6.162010000e-07 V_low
+ 6.163000000e-07 V_low
+ 6.163010000e-07 V_low
+ 6.164000000e-07 V_low
+ 6.164010000e-07 V_low
+ 6.165000000e-07 V_low
+ 6.165010000e-07 V_low
+ 6.166000000e-07 V_low
+ 6.166010000e-07 V_low
+ 6.167000000e-07 V_low
+ 6.167010000e-07 V_low
+ 6.168000000e-07 V_low
+ 6.168010000e-07 V_low
+ 6.169000000e-07 V_low
+ 6.169010000e-07 V_hig
+ 6.170000000e-07 V_hig
+ 6.170010000e-07 V_hig
+ 6.171000000e-07 V_hig
+ 6.171010000e-07 V_hig
+ 6.172000000e-07 V_hig
+ 6.172010000e-07 V_hig
+ 6.173000000e-07 V_hig
+ 6.173010000e-07 V_hig
+ 6.174000000e-07 V_hig
+ 6.174010000e-07 V_hig
+ 6.175000000e-07 V_hig
+ 6.175010000e-07 V_hig
+ 6.176000000e-07 V_hig
+ 6.176010000e-07 V_hig
+ 6.177000000e-07 V_hig
+ 6.177010000e-07 V_hig
+ 6.178000000e-07 V_hig
+ 6.178010000e-07 V_hig
+ 6.179000000e-07 V_hig
+ 6.179010000e-07 V_hig
+ 6.180000000e-07 V_hig
+ 6.180010000e-07 V_hig
+ 6.181000000e-07 V_hig
+ 6.181010000e-07 V_hig
+ 6.182000000e-07 V_hig
+ 6.182010000e-07 V_hig
+ 6.183000000e-07 V_hig
+ 6.183010000e-07 V_hig
+ 6.184000000e-07 V_hig
+ 6.184010000e-07 V_hig
+ 6.185000000e-07 V_hig
+ 6.185010000e-07 V_hig
+ 6.186000000e-07 V_hig
+ 6.186010000e-07 V_hig
+ 6.187000000e-07 V_hig
+ 6.187010000e-07 V_hig
+ 6.188000000e-07 V_hig
+ 6.188010000e-07 V_hig
+ 6.189000000e-07 V_hig
+ 6.189010000e-07 V_low
+ 6.190000000e-07 V_low
+ 6.190010000e-07 V_low
+ 6.191000000e-07 V_low
+ 6.191010000e-07 V_low
+ 6.192000000e-07 V_low
+ 6.192010000e-07 V_low
+ 6.193000000e-07 V_low
+ 6.193010000e-07 V_low
+ 6.194000000e-07 V_low
+ 6.194010000e-07 V_low
+ 6.195000000e-07 V_low
+ 6.195010000e-07 V_low
+ 6.196000000e-07 V_low
+ 6.196010000e-07 V_low
+ 6.197000000e-07 V_low
+ 6.197010000e-07 V_low
+ 6.198000000e-07 V_low
+ 6.198010000e-07 V_low
+ 6.199000000e-07 V_low
+ 6.199010000e-07 V_low
+ 6.200000000e-07 V_low
+ 6.200010000e-07 V_low
+ 6.201000000e-07 V_low
+ 6.201010000e-07 V_low
+ 6.202000000e-07 V_low
+ 6.202010000e-07 V_low
+ 6.203000000e-07 V_low
+ 6.203010000e-07 V_low
+ 6.204000000e-07 V_low
+ 6.204010000e-07 V_low
+ 6.205000000e-07 V_low
+ 6.205010000e-07 V_low
+ 6.206000000e-07 V_low
+ 6.206010000e-07 V_low
+ 6.207000000e-07 V_low
+ 6.207010000e-07 V_low
+ 6.208000000e-07 V_low
+ 6.208010000e-07 V_low
+ 6.209000000e-07 V_low
+ 6.209010000e-07 V_hig
+ 6.210000000e-07 V_hig
+ 6.210010000e-07 V_hig
+ 6.211000000e-07 V_hig
+ 6.211010000e-07 V_hig
+ 6.212000000e-07 V_hig
+ 6.212010000e-07 V_hig
+ 6.213000000e-07 V_hig
+ 6.213010000e-07 V_hig
+ 6.214000000e-07 V_hig
+ 6.214010000e-07 V_hig
+ 6.215000000e-07 V_hig
+ 6.215010000e-07 V_hig
+ 6.216000000e-07 V_hig
+ 6.216010000e-07 V_hig
+ 6.217000000e-07 V_hig
+ 6.217010000e-07 V_hig
+ 6.218000000e-07 V_hig
+ 6.218010000e-07 V_hig
+ 6.219000000e-07 V_hig
+ 6.219010000e-07 V_hig
+ 6.220000000e-07 V_hig
+ 6.220010000e-07 V_hig
+ 6.221000000e-07 V_hig
+ 6.221010000e-07 V_hig
+ 6.222000000e-07 V_hig
+ 6.222010000e-07 V_hig
+ 6.223000000e-07 V_hig
+ 6.223010000e-07 V_hig
+ 6.224000000e-07 V_hig
+ 6.224010000e-07 V_hig
+ 6.225000000e-07 V_hig
+ 6.225010000e-07 V_hig
+ 6.226000000e-07 V_hig
+ 6.226010000e-07 V_hig
+ 6.227000000e-07 V_hig
+ 6.227010000e-07 V_hig
+ 6.228000000e-07 V_hig
+ 6.228010000e-07 V_hig
+ 6.229000000e-07 V_hig
+ 6.229010000e-07 V_low
+ 6.230000000e-07 V_low
+ 6.230010000e-07 V_low
+ 6.231000000e-07 V_low
+ 6.231010000e-07 V_low
+ 6.232000000e-07 V_low
+ 6.232010000e-07 V_low
+ 6.233000000e-07 V_low
+ 6.233010000e-07 V_low
+ 6.234000000e-07 V_low
+ 6.234010000e-07 V_low
+ 6.235000000e-07 V_low
+ 6.235010000e-07 V_low
+ 6.236000000e-07 V_low
+ 6.236010000e-07 V_low
+ 6.237000000e-07 V_low
+ 6.237010000e-07 V_low
+ 6.238000000e-07 V_low
+ 6.238010000e-07 V_low
+ 6.239000000e-07 V_low
+ 6.239010000e-07 V_hig
+ 6.240000000e-07 V_hig
+ 6.240010000e-07 V_hig
+ 6.241000000e-07 V_hig
+ 6.241010000e-07 V_hig
+ 6.242000000e-07 V_hig
+ 6.242010000e-07 V_hig
+ 6.243000000e-07 V_hig
+ 6.243010000e-07 V_hig
+ 6.244000000e-07 V_hig
+ 6.244010000e-07 V_hig
+ 6.245000000e-07 V_hig
+ 6.245010000e-07 V_hig
+ 6.246000000e-07 V_hig
+ 6.246010000e-07 V_hig
+ 6.247000000e-07 V_hig
+ 6.247010000e-07 V_hig
+ 6.248000000e-07 V_hig
+ 6.248010000e-07 V_hig
+ 6.249000000e-07 V_hig
+ 6.249010000e-07 V_low
+ 6.250000000e-07 V_low
+ 6.250010000e-07 V_low
+ 6.251000000e-07 V_low
+ 6.251010000e-07 V_low
+ 6.252000000e-07 V_low
+ 6.252010000e-07 V_low
+ 6.253000000e-07 V_low
+ 6.253010000e-07 V_low
+ 6.254000000e-07 V_low
+ 6.254010000e-07 V_low
+ 6.255000000e-07 V_low
+ 6.255010000e-07 V_low
+ 6.256000000e-07 V_low
+ 6.256010000e-07 V_low
+ 6.257000000e-07 V_low
+ 6.257010000e-07 V_low
+ 6.258000000e-07 V_low
+ 6.258010000e-07 V_low
+ 6.259000000e-07 V_low
+ 6.259010000e-07 V_low
+ 6.260000000e-07 V_low
+ 6.260010000e-07 V_low
+ 6.261000000e-07 V_low
+ 6.261010000e-07 V_low
+ 6.262000000e-07 V_low
+ 6.262010000e-07 V_low
+ 6.263000000e-07 V_low
+ 6.263010000e-07 V_low
+ 6.264000000e-07 V_low
+ 6.264010000e-07 V_low
+ 6.265000000e-07 V_low
+ 6.265010000e-07 V_low
+ 6.266000000e-07 V_low
+ 6.266010000e-07 V_low
+ 6.267000000e-07 V_low
+ 6.267010000e-07 V_low
+ 6.268000000e-07 V_low
+ 6.268010000e-07 V_low
+ 6.269000000e-07 V_low
+ 6.269010000e-07 V_low
+ 6.270000000e-07 V_low
+ 6.270010000e-07 V_low
+ 6.271000000e-07 V_low
+ 6.271010000e-07 V_low
+ 6.272000000e-07 V_low
+ 6.272010000e-07 V_low
+ 6.273000000e-07 V_low
+ 6.273010000e-07 V_low
+ 6.274000000e-07 V_low
+ 6.274010000e-07 V_low
+ 6.275000000e-07 V_low
+ 6.275010000e-07 V_low
+ 6.276000000e-07 V_low
+ 6.276010000e-07 V_low
+ 6.277000000e-07 V_low
+ 6.277010000e-07 V_low
+ 6.278000000e-07 V_low
+ 6.278010000e-07 V_low
+ 6.279000000e-07 V_low
+ 6.279010000e-07 V_hig
+ 6.280000000e-07 V_hig
+ 6.280010000e-07 V_hig
+ 6.281000000e-07 V_hig
+ 6.281010000e-07 V_hig
+ 6.282000000e-07 V_hig
+ 6.282010000e-07 V_hig
+ 6.283000000e-07 V_hig
+ 6.283010000e-07 V_hig
+ 6.284000000e-07 V_hig
+ 6.284010000e-07 V_hig
+ 6.285000000e-07 V_hig
+ 6.285010000e-07 V_hig
+ 6.286000000e-07 V_hig
+ 6.286010000e-07 V_hig
+ 6.287000000e-07 V_hig
+ 6.287010000e-07 V_hig
+ 6.288000000e-07 V_hig
+ 6.288010000e-07 V_hig
+ 6.289000000e-07 V_hig
+ 6.289010000e-07 V_hig
+ 6.290000000e-07 V_hig
+ 6.290010000e-07 V_hig
+ 6.291000000e-07 V_hig
+ 6.291010000e-07 V_hig
+ 6.292000000e-07 V_hig
+ 6.292010000e-07 V_hig
+ 6.293000000e-07 V_hig
+ 6.293010000e-07 V_hig
+ 6.294000000e-07 V_hig
+ 6.294010000e-07 V_hig
+ 6.295000000e-07 V_hig
+ 6.295010000e-07 V_hig
+ 6.296000000e-07 V_hig
+ 6.296010000e-07 V_hig
+ 6.297000000e-07 V_hig
+ 6.297010000e-07 V_hig
+ 6.298000000e-07 V_hig
+ 6.298010000e-07 V_hig
+ 6.299000000e-07 V_hig
+ 6.299010000e-07 V_hig
+ 6.300000000e-07 V_hig
+ 6.300010000e-07 V_hig
+ 6.301000000e-07 V_hig
+ 6.301010000e-07 V_hig
+ 6.302000000e-07 V_hig
+ 6.302010000e-07 V_hig
+ 6.303000000e-07 V_hig
+ 6.303010000e-07 V_hig
+ 6.304000000e-07 V_hig
+ 6.304010000e-07 V_hig
+ 6.305000000e-07 V_hig
+ 6.305010000e-07 V_hig
+ 6.306000000e-07 V_hig
+ 6.306010000e-07 V_hig
+ 6.307000000e-07 V_hig
+ 6.307010000e-07 V_hig
+ 6.308000000e-07 V_hig
+ 6.308010000e-07 V_hig
+ 6.309000000e-07 V_hig
+ 6.309010000e-07 V_hig
+ 6.310000000e-07 V_hig
+ 6.310010000e-07 V_hig
+ 6.311000000e-07 V_hig
+ 6.311010000e-07 V_hig
+ 6.312000000e-07 V_hig
+ 6.312010000e-07 V_hig
+ 6.313000000e-07 V_hig
+ 6.313010000e-07 V_hig
+ 6.314000000e-07 V_hig
+ 6.314010000e-07 V_hig
+ 6.315000000e-07 V_hig
+ 6.315010000e-07 V_hig
+ 6.316000000e-07 V_hig
+ 6.316010000e-07 V_hig
+ 6.317000000e-07 V_hig
+ 6.317010000e-07 V_hig
+ 6.318000000e-07 V_hig
+ 6.318010000e-07 V_hig
+ 6.319000000e-07 V_hig
+ 6.319010000e-07 V_low
+ 6.320000000e-07 V_low
+ 6.320010000e-07 V_low
+ 6.321000000e-07 V_low
+ 6.321010000e-07 V_low
+ 6.322000000e-07 V_low
+ 6.322010000e-07 V_low
+ 6.323000000e-07 V_low
+ 6.323010000e-07 V_low
+ 6.324000000e-07 V_low
+ 6.324010000e-07 V_low
+ 6.325000000e-07 V_low
+ 6.325010000e-07 V_low
+ 6.326000000e-07 V_low
+ 6.326010000e-07 V_low
+ 6.327000000e-07 V_low
+ 6.327010000e-07 V_low
+ 6.328000000e-07 V_low
+ 6.328010000e-07 V_low
+ 6.329000000e-07 V_low
+ 6.329010000e-07 V_low
+ 6.330000000e-07 V_low
+ 6.330010000e-07 V_low
+ 6.331000000e-07 V_low
+ 6.331010000e-07 V_low
+ 6.332000000e-07 V_low
+ 6.332010000e-07 V_low
+ 6.333000000e-07 V_low
+ 6.333010000e-07 V_low
+ 6.334000000e-07 V_low
+ 6.334010000e-07 V_low
+ 6.335000000e-07 V_low
+ 6.335010000e-07 V_low
+ 6.336000000e-07 V_low
+ 6.336010000e-07 V_low
+ 6.337000000e-07 V_low
+ 6.337010000e-07 V_low
+ 6.338000000e-07 V_low
+ 6.338010000e-07 V_low
+ 6.339000000e-07 V_low
+ 6.339010000e-07 V_hig
+ 6.340000000e-07 V_hig
+ 6.340010000e-07 V_hig
+ 6.341000000e-07 V_hig
+ 6.341010000e-07 V_hig
+ 6.342000000e-07 V_hig
+ 6.342010000e-07 V_hig
+ 6.343000000e-07 V_hig
+ 6.343010000e-07 V_hig
+ 6.344000000e-07 V_hig
+ 6.344010000e-07 V_hig
+ 6.345000000e-07 V_hig
+ 6.345010000e-07 V_hig
+ 6.346000000e-07 V_hig
+ 6.346010000e-07 V_hig
+ 6.347000000e-07 V_hig
+ 6.347010000e-07 V_hig
+ 6.348000000e-07 V_hig
+ 6.348010000e-07 V_hig
+ 6.349000000e-07 V_hig
+ 6.349010000e-07 V_low
+ 6.350000000e-07 V_low
+ 6.350010000e-07 V_low
+ 6.351000000e-07 V_low
+ 6.351010000e-07 V_low
+ 6.352000000e-07 V_low
+ 6.352010000e-07 V_low
+ 6.353000000e-07 V_low
+ 6.353010000e-07 V_low
+ 6.354000000e-07 V_low
+ 6.354010000e-07 V_low
+ 6.355000000e-07 V_low
+ 6.355010000e-07 V_low
+ 6.356000000e-07 V_low
+ 6.356010000e-07 V_low
+ 6.357000000e-07 V_low
+ 6.357010000e-07 V_low
+ 6.358000000e-07 V_low
+ 6.358010000e-07 V_low
+ 6.359000000e-07 V_low
+ 6.359010000e-07 V_hig
+ 6.360000000e-07 V_hig
+ 6.360010000e-07 V_hig
+ 6.361000000e-07 V_hig
+ 6.361010000e-07 V_hig
+ 6.362000000e-07 V_hig
+ 6.362010000e-07 V_hig
+ 6.363000000e-07 V_hig
+ 6.363010000e-07 V_hig
+ 6.364000000e-07 V_hig
+ 6.364010000e-07 V_hig
+ 6.365000000e-07 V_hig
+ 6.365010000e-07 V_hig
+ 6.366000000e-07 V_hig
+ 6.366010000e-07 V_hig
+ 6.367000000e-07 V_hig
+ 6.367010000e-07 V_hig
+ 6.368000000e-07 V_hig
+ 6.368010000e-07 V_hig
+ 6.369000000e-07 V_hig
+ 6.369010000e-07 V_hig
+ 6.370000000e-07 V_hig
+ 6.370010000e-07 V_hig
+ 6.371000000e-07 V_hig
+ 6.371010000e-07 V_hig
+ 6.372000000e-07 V_hig
+ 6.372010000e-07 V_hig
+ 6.373000000e-07 V_hig
+ 6.373010000e-07 V_hig
+ 6.374000000e-07 V_hig
+ 6.374010000e-07 V_hig
+ 6.375000000e-07 V_hig
+ 6.375010000e-07 V_hig
+ 6.376000000e-07 V_hig
+ 6.376010000e-07 V_hig
+ 6.377000000e-07 V_hig
+ 6.377010000e-07 V_hig
+ 6.378000000e-07 V_hig
+ 6.378010000e-07 V_hig
+ 6.379000000e-07 V_hig
+ 6.379010000e-07 V_hig
+ 6.380000000e-07 V_hig
+ 6.380010000e-07 V_hig
+ 6.381000000e-07 V_hig
+ 6.381010000e-07 V_hig
+ 6.382000000e-07 V_hig
+ 6.382010000e-07 V_hig
+ 6.383000000e-07 V_hig
+ 6.383010000e-07 V_hig
+ 6.384000000e-07 V_hig
+ 6.384010000e-07 V_hig
+ 6.385000000e-07 V_hig
+ 6.385010000e-07 V_hig
+ 6.386000000e-07 V_hig
+ 6.386010000e-07 V_hig
+ 6.387000000e-07 V_hig
+ 6.387010000e-07 V_hig
+ 6.388000000e-07 V_hig
+ 6.388010000e-07 V_hig
+ 6.389000000e-07 V_hig
+ 6.389010000e-07 V_low
+ 6.390000000e-07 V_low
+ 6.390010000e-07 V_low
+ 6.391000000e-07 V_low
+ 6.391010000e-07 V_low
+ 6.392000000e-07 V_low
+ 6.392010000e-07 V_low
+ 6.393000000e-07 V_low
+ 6.393010000e-07 V_low
+ 6.394000000e-07 V_low
+ 6.394010000e-07 V_low
+ 6.395000000e-07 V_low
+ 6.395010000e-07 V_low
+ 6.396000000e-07 V_low
+ 6.396010000e-07 V_low
+ 6.397000000e-07 V_low
+ 6.397010000e-07 V_low
+ 6.398000000e-07 V_low
+ 6.398010000e-07 V_low
+ 6.399000000e-07 V_low
+ 6.399010000e-07 V_hig
+ 6.400000000e-07 V_hig
+ 6.400010000e-07 V_hig
+ 6.401000000e-07 V_hig
+ 6.401010000e-07 V_hig
+ 6.402000000e-07 V_hig
+ 6.402010000e-07 V_hig
+ 6.403000000e-07 V_hig
+ 6.403010000e-07 V_hig
+ 6.404000000e-07 V_hig
+ 6.404010000e-07 V_hig
+ 6.405000000e-07 V_hig
+ 6.405010000e-07 V_hig
+ 6.406000000e-07 V_hig
+ 6.406010000e-07 V_hig
+ 6.407000000e-07 V_hig
+ 6.407010000e-07 V_hig
+ 6.408000000e-07 V_hig
+ 6.408010000e-07 V_hig
+ 6.409000000e-07 V_hig
+ 6.409010000e-07 V_hig
+ 6.410000000e-07 V_hig
+ 6.410010000e-07 V_hig
+ 6.411000000e-07 V_hig
+ 6.411010000e-07 V_hig
+ 6.412000000e-07 V_hig
+ 6.412010000e-07 V_hig
+ 6.413000000e-07 V_hig
+ 6.413010000e-07 V_hig
+ 6.414000000e-07 V_hig
+ 6.414010000e-07 V_hig
+ 6.415000000e-07 V_hig
+ 6.415010000e-07 V_hig
+ 6.416000000e-07 V_hig
+ 6.416010000e-07 V_hig
+ 6.417000000e-07 V_hig
+ 6.417010000e-07 V_hig
+ 6.418000000e-07 V_hig
+ 6.418010000e-07 V_hig
+ 6.419000000e-07 V_hig
+ 6.419010000e-07 V_hig
+ 6.420000000e-07 V_hig
+ 6.420010000e-07 V_hig
+ 6.421000000e-07 V_hig
+ 6.421010000e-07 V_hig
+ 6.422000000e-07 V_hig
+ 6.422010000e-07 V_hig
+ 6.423000000e-07 V_hig
+ 6.423010000e-07 V_hig
+ 6.424000000e-07 V_hig
+ 6.424010000e-07 V_hig
+ 6.425000000e-07 V_hig
+ 6.425010000e-07 V_hig
+ 6.426000000e-07 V_hig
+ 6.426010000e-07 V_hig
+ 6.427000000e-07 V_hig
+ 6.427010000e-07 V_hig
+ 6.428000000e-07 V_hig
+ 6.428010000e-07 V_hig
+ 6.429000000e-07 V_hig
+ 6.429010000e-07 V_hig
+ 6.430000000e-07 V_hig
+ 6.430010000e-07 V_hig
+ 6.431000000e-07 V_hig
+ 6.431010000e-07 V_hig
+ 6.432000000e-07 V_hig
+ 6.432010000e-07 V_hig
+ 6.433000000e-07 V_hig
+ 6.433010000e-07 V_hig
+ 6.434000000e-07 V_hig
+ 6.434010000e-07 V_hig
+ 6.435000000e-07 V_hig
+ 6.435010000e-07 V_hig
+ 6.436000000e-07 V_hig
+ 6.436010000e-07 V_hig
+ 6.437000000e-07 V_hig
+ 6.437010000e-07 V_hig
+ 6.438000000e-07 V_hig
+ 6.438010000e-07 V_hig
+ 6.439000000e-07 V_hig
+ 6.439010000e-07 V_hig
+ 6.440000000e-07 V_hig
+ 6.440010000e-07 V_hig
+ 6.441000000e-07 V_hig
+ 6.441010000e-07 V_hig
+ 6.442000000e-07 V_hig
+ 6.442010000e-07 V_hig
+ 6.443000000e-07 V_hig
+ 6.443010000e-07 V_hig
+ 6.444000000e-07 V_hig
+ 6.444010000e-07 V_hig
+ 6.445000000e-07 V_hig
+ 6.445010000e-07 V_hig
+ 6.446000000e-07 V_hig
+ 6.446010000e-07 V_hig
+ 6.447000000e-07 V_hig
+ 6.447010000e-07 V_hig
+ 6.448000000e-07 V_hig
+ 6.448010000e-07 V_hig
+ 6.449000000e-07 V_hig
+ 6.449010000e-07 V_low
+ 6.450000000e-07 V_low
+ 6.450010000e-07 V_low
+ 6.451000000e-07 V_low
+ 6.451010000e-07 V_low
+ 6.452000000e-07 V_low
+ 6.452010000e-07 V_low
+ 6.453000000e-07 V_low
+ 6.453010000e-07 V_low
+ 6.454000000e-07 V_low
+ 6.454010000e-07 V_low
+ 6.455000000e-07 V_low
+ 6.455010000e-07 V_low
+ 6.456000000e-07 V_low
+ 6.456010000e-07 V_low
+ 6.457000000e-07 V_low
+ 6.457010000e-07 V_low
+ 6.458000000e-07 V_low
+ 6.458010000e-07 V_low
+ 6.459000000e-07 V_low
+ 6.459010000e-07 V_hig
+ 6.460000000e-07 V_hig
+ 6.460010000e-07 V_hig
+ 6.461000000e-07 V_hig
+ 6.461010000e-07 V_hig
+ 6.462000000e-07 V_hig
+ 6.462010000e-07 V_hig
+ 6.463000000e-07 V_hig
+ 6.463010000e-07 V_hig
+ 6.464000000e-07 V_hig
+ 6.464010000e-07 V_hig
+ 6.465000000e-07 V_hig
+ 6.465010000e-07 V_hig
+ 6.466000000e-07 V_hig
+ 6.466010000e-07 V_hig
+ 6.467000000e-07 V_hig
+ 6.467010000e-07 V_hig
+ 6.468000000e-07 V_hig
+ 6.468010000e-07 V_hig
+ 6.469000000e-07 V_hig
+ 6.469010000e-07 V_hig
+ 6.470000000e-07 V_hig
+ 6.470010000e-07 V_hig
+ 6.471000000e-07 V_hig
+ 6.471010000e-07 V_hig
+ 6.472000000e-07 V_hig
+ 6.472010000e-07 V_hig
+ 6.473000000e-07 V_hig
+ 6.473010000e-07 V_hig
+ 6.474000000e-07 V_hig
+ 6.474010000e-07 V_hig
+ 6.475000000e-07 V_hig
+ 6.475010000e-07 V_hig
+ 6.476000000e-07 V_hig
+ 6.476010000e-07 V_hig
+ 6.477000000e-07 V_hig
+ 6.477010000e-07 V_hig
+ 6.478000000e-07 V_hig
+ 6.478010000e-07 V_hig
+ 6.479000000e-07 V_hig
+ 6.479010000e-07 V_hig
+ 6.480000000e-07 V_hig
+ 6.480010000e-07 V_hig
+ 6.481000000e-07 V_hig
+ 6.481010000e-07 V_hig
+ 6.482000000e-07 V_hig
+ 6.482010000e-07 V_hig
+ 6.483000000e-07 V_hig
+ 6.483010000e-07 V_hig
+ 6.484000000e-07 V_hig
+ 6.484010000e-07 V_hig
+ 6.485000000e-07 V_hig
+ 6.485010000e-07 V_hig
+ 6.486000000e-07 V_hig
+ 6.486010000e-07 V_hig
+ 6.487000000e-07 V_hig
+ 6.487010000e-07 V_hig
+ 6.488000000e-07 V_hig
+ 6.488010000e-07 V_hig
+ 6.489000000e-07 V_hig
+ 6.489010000e-07 V_low
+ 6.490000000e-07 V_low
+ 6.490010000e-07 V_low
+ 6.491000000e-07 V_low
+ 6.491010000e-07 V_low
+ 6.492000000e-07 V_low
+ 6.492010000e-07 V_low
+ 6.493000000e-07 V_low
+ 6.493010000e-07 V_low
+ 6.494000000e-07 V_low
+ 6.494010000e-07 V_low
+ 6.495000000e-07 V_low
+ 6.495010000e-07 V_low
+ 6.496000000e-07 V_low
+ 6.496010000e-07 V_low
+ 6.497000000e-07 V_low
+ 6.497010000e-07 V_low
+ 6.498000000e-07 V_low
+ 6.498010000e-07 V_low
+ 6.499000000e-07 V_low
+ 6.499010000e-07 V_hig
+ 6.500000000e-07 V_hig
+ 6.500010000e-07 V_hig
+ 6.501000000e-07 V_hig
+ 6.501010000e-07 V_hig
+ 6.502000000e-07 V_hig
+ 6.502010000e-07 V_hig
+ 6.503000000e-07 V_hig
+ 6.503010000e-07 V_hig
+ 6.504000000e-07 V_hig
+ 6.504010000e-07 V_hig
+ 6.505000000e-07 V_hig
+ 6.505010000e-07 V_hig
+ 6.506000000e-07 V_hig
+ 6.506010000e-07 V_hig
+ 6.507000000e-07 V_hig
+ 6.507010000e-07 V_hig
+ 6.508000000e-07 V_hig
+ 6.508010000e-07 V_hig
+ 6.509000000e-07 V_hig
+ 6.509010000e-07 V_hig
+ 6.510000000e-07 V_hig
+ 6.510010000e-07 V_hig
+ 6.511000000e-07 V_hig
+ 6.511010000e-07 V_hig
+ 6.512000000e-07 V_hig
+ 6.512010000e-07 V_hig
+ 6.513000000e-07 V_hig
+ 6.513010000e-07 V_hig
+ 6.514000000e-07 V_hig
+ 6.514010000e-07 V_hig
+ 6.515000000e-07 V_hig
+ 6.515010000e-07 V_hig
+ 6.516000000e-07 V_hig
+ 6.516010000e-07 V_hig
+ 6.517000000e-07 V_hig
+ 6.517010000e-07 V_hig
+ 6.518000000e-07 V_hig
+ 6.518010000e-07 V_hig
+ 6.519000000e-07 V_hig
+ 6.519010000e-07 V_hig
+ 6.520000000e-07 V_hig
+ 6.520010000e-07 V_hig
+ 6.521000000e-07 V_hig
+ 6.521010000e-07 V_hig
+ 6.522000000e-07 V_hig
+ 6.522010000e-07 V_hig
+ 6.523000000e-07 V_hig
+ 6.523010000e-07 V_hig
+ 6.524000000e-07 V_hig
+ 6.524010000e-07 V_hig
+ 6.525000000e-07 V_hig
+ 6.525010000e-07 V_hig
+ 6.526000000e-07 V_hig
+ 6.526010000e-07 V_hig
+ 6.527000000e-07 V_hig
+ 6.527010000e-07 V_hig
+ 6.528000000e-07 V_hig
+ 6.528010000e-07 V_hig
+ 6.529000000e-07 V_hig
+ 6.529010000e-07 V_hig
+ 6.530000000e-07 V_hig
+ 6.530010000e-07 V_hig
+ 6.531000000e-07 V_hig
+ 6.531010000e-07 V_hig
+ 6.532000000e-07 V_hig
+ 6.532010000e-07 V_hig
+ 6.533000000e-07 V_hig
+ 6.533010000e-07 V_hig
+ 6.534000000e-07 V_hig
+ 6.534010000e-07 V_hig
+ 6.535000000e-07 V_hig
+ 6.535010000e-07 V_hig
+ 6.536000000e-07 V_hig
+ 6.536010000e-07 V_hig
+ 6.537000000e-07 V_hig
+ 6.537010000e-07 V_hig
+ 6.538000000e-07 V_hig
+ 6.538010000e-07 V_hig
+ 6.539000000e-07 V_hig
+ 6.539010000e-07 V_low
+ 6.540000000e-07 V_low
+ 6.540010000e-07 V_low
+ 6.541000000e-07 V_low
+ 6.541010000e-07 V_low
+ 6.542000000e-07 V_low
+ 6.542010000e-07 V_low
+ 6.543000000e-07 V_low
+ 6.543010000e-07 V_low
+ 6.544000000e-07 V_low
+ 6.544010000e-07 V_low
+ 6.545000000e-07 V_low
+ 6.545010000e-07 V_low
+ 6.546000000e-07 V_low
+ 6.546010000e-07 V_low
+ 6.547000000e-07 V_low
+ 6.547010000e-07 V_low
+ 6.548000000e-07 V_low
+ 6.548010000e-07 V_low
+ 6.549000000e-07 V_low
+ 6.549010000e-07 V_low
+ 6.550000000e-07 V_low
+ 6.550010000e-07 V_low
+ 6.551000000e-07 V_low
+ 6.551010000e-07 V_low
+ 6.552000000e-07 V_low
+ 6.552010000e-07 V_low
+ 6.553000000e-07 V_low
+ 6.553010000e-07 V_low
+ 6.554000000e-07 V_low
+ 6.554010000e-07 V_low
+ 6.555000000e-07 V_low
+ 6.555010000e-07 V_low
+ 6.556000000e-07 V_low
+ 6.556010000e-07 V_low
+ 6.557000000e-07 V_low
+ 6.557010000e-07 V_low
+ 6.558000000e-07 V_low
+ 6.558010000e-07 V_low
+ 6.559000000e-07 V_low
+ 6.559010000e-07 V_hig
+ 6.560000000e-07 V_hig
+ 6.560010000e-07 V_hig
+ 6.561000000e-07 V_hig
+ 6.561010000e-07 V_hig
+ 6.562000000e-07 V_hig
+ 6.562010000e-07 V_hig
+ 6.563000000e-07 V_hig
+ 6.563010000e-07 V_hig
+ 6.564000000e-07 V_hig
+ 6.564010000e-07 V_hig
+ 6.565000000e-07 V_hig
+ 6.565010000e-07 V_hig
+ 6.566000000e-07 V_hig
+ 6.566010000e-07 V_hig
+ 6.567000000e-07 V_hig
+ 6.567010000e-07 V_hig
+ 6.568000000e-07 V_hig
+ 6.568010000e-07 V_hig
+ 6.569000000e-07 V_hig
+ 6.569010000e-07 V_low
+ 6.570000000e-07 V_low
+ 6.570010000e-07 V_low
+ 6.571000000e-07 V_low
+ 6.571010000e-07 V_low
+ 6.572000000e-07 V_low
+ 6.572010000e-07 V_low
+ 6.573000000e-07 V_low
+ 6.573010000e-07 V_low
+ 6.574000000e-07 V_low
+ 6.574010000e-07 V_low
+ 6.575000000e-07 V_low
+ 6.575010000e-07 V_low
+ 6.576000000e-07 V_low
+ 6.576010000e-07 V_low
+ 6.577000000e-07 V_low
+ 6.577010000e-07 V_low
+ 6.578000000e-07 V_low
+ 6.578010000e-07 V_low
+ 6.579000000e-07 V_low
+ 6.579010000e-07 V_low
+ 6.580000000e-07 V_low
+ 6.580010000e-07 V_low
+ 6.581000000e-07 V_low
+ 6.581010000e-07 V_low
+ 6.582000000e-07 V_low
+ 6.582010000e-07 V_low
+ 6.583000000e-07 V_low
+ 6.583010000e-07 V_low
+ 6.584000000e-07 V_low
+ 6.584010000e-07 V_low
+ 6.585000000e-07 V_low
+ 6.585010000e-07 V_low
+ 6.586000000e-07 V_low
+ 6.586010000e-07 V_low
+ 6.587000000e-07 V_low
+ 6.587010000e-07 V_low
+ 6.588000000e-07 V_low
+ 6.588010000e-07 V_low
+ 6.589000000e-07 V_low
+ 6.589010000e-07 V_hig
+ 6.590000000e-07 V_hig
+ 6.590010000e-07 V_hig
+ 6.591000000e-07 V_hig
+ 6.591010000e-07 V_hig
+ 6.592000000e-07 V_hig
+ 6.592010000e-07 V_hig
+ 6.593000000e-07 V_hig
+ 6.593010000e-07 V_hig
+ 6.594000000e-07 V_hig
+ 6.594010000e-07 V_hig
+ 6.595000000e-07 V_hig
+ 6.595010000e-07 V_hig
+ 6.596000000e-07 V_hig
+ 6.596010000e-07 V_hig
+ 6.597000000e-07 V_hig
+ 6.597010000e-07 V_hig
+ 6.598000000e-07 V_hig
+ 6.598010000e-07 V_hig
+ 6.599000000e-07 V_hig
+ 6.599010000e-07 V_low
+ 6.600000000e-07 V_low
+ 6.600010000e-07 V_low
+ 6.601000000e-07 V_low
+ 6.601010000e-07 V_low
+ 6.602000000e-07 V_low
+ 6.602010000e-07 V_low
+ 6.603000000e-07 V_low
+ 6.603010000e-07 V_low
+ 6.604000000e-07 V_low
+ 6.604010000e-07 V_low
+ 6.605000000e-07 V_low
+ 6.605010000e-07 V_low
+ 6.606000000e-07 V_low
+ 6.606010000e-07 V_low
+ 6.607000000e-07 V_low
+ 6.607010000e-07 V_low
+ 6.608000000e-07 V_low
+ 6.608010000e-07 V_low
+ 6.609000000e-07 V_low
+ 6.609010000e-07 V_hig
+ 6.610000000e-07 V_hig
+ 6.610010000e-07 V_hig
+ 6.611000000e-07 V_hig
+ 6.611010000e-07 V_hig
+ 6.612000000e-07 V_hig
+ 6.612010000e-07 V_hig
+ 6.613000000e-07 V_hig
+ 6.613010000e-07 V_hig
+ 6.614000000e-07 V_hig
+ 6.614010000e-07 V_hig
+ 6.615000000e-07 V_hig
+ 6.615010000e-07 V_hig
+ 6.616000000e-07 V_hig
+ 6.616010000e-07 V_hig
+ 6.617000000e-07 V_hig
+ 6.617010000e-07 V_hig
+ 6.618000000e-07 V_hig
+ 6.618010000e-07 V_hig
+ 6.619000000e-07 V_hig
+ 6.619010000e-07 V_hig
+ 6.620000000e-07 V_hig
+ 6.620010000e-07 V_hig
+ 6.621000000e-07 V_hig
+ 6.621010000e-07 V_hig
+ 6.622000000e-07 V_hig
+ 6.622010000e-07 V_hig
+ 6.623000000e-07 V_hig
+ 6.623010000e-07 V_hig
+ 6.624000000e-07 V_hig
+ 6.624010000e-07 V_hig
+ 6.625000000e-07 V_hig
+ 6.625010000e-07 V_hig
+ 6.626000000e-07 V_hig
+ 6.626010000e-07 V_hig
+ 6.627000000e-07 V_hig
+ 6.627010000e-07 V_hig
+ 6.628000000e-07 V_hig
+ 6.628010000e-07 V_hig
+ 6.629000000e-07 V_hig
+ 6.629010000e-07 V_hig
+ 6.630000000e-07 V_hig
+ 6.630010000e-07 V_hig
+ 6.631000000e-07 V_hig
+ 6.631010000e-07 V_hig
+ 6.632000000e-07 V_hig
+ 6.632010000e-07 V_hig
+ 6.633000000e-07 V_hig
+ 6.633010000e-07 V_hig
+ 6.634000000e-07 V_hig
+ 6.634010000e-07 V_hig
+ 6.635000000e-07 V_hig
+ 6.635010000e-07 V_hig
+ 6.636000000e-07 V_hig
+ 6.636010000e-07 V_hig
+ 6.637000000e-07 V_hig
+ 6.637010000e-07 V_hig
+ 6.638000000e-07 V_hig
+ 6.638010000e-07 V_hig
+ 6.639000000e-07 V_hig
+ 6.639010000e-07 V_hig
+ 6.640000000e-07 V_hig
+ 6.640010000e-07 V_hig
+ 6.641000000e-07 V_hig
+ 6.641010000e-07 V_hig
+ 6.642000000e-07 V_hig
+ 6.642010000e-07 V_hig
+ 6.643000000e-07 V_hig
+ 6.643010000e-07 V_hig
+ 6.644000000e-07 V_hig
+ 6.644010000e-07 V_hig
+ 6.645000000e-07 V_hig
+ 6.645010000e-07 V_hig
+ 6.646000000e-07 V_hig
+ 6.646010000e-07 V_hig
+ 6.647000000e-07 V_hig
+ 6.647010000e-07 V_hig
+ 6.648000000e-07 V_hig
+ 6.648010000e-07 V_hig
+ 6.649000000e-07 V_hig
+ 6.649010000e-07 V_hig
+ 6.650000000e-07 V_hig
+ 6.650010000e-07 V_hig
+ 6.651000000e-07 V_hig
+ 6.651010000e-07 V_hig
+ 6.652000000e-07 V_hig
+ 6.652010000e-07 V_hig
+ 6.653000000e-07 V_hig
+ 6.653010000e-07 V_hig
+ 6.654000000e-07 V_hig
+ 6.654010000e-07 V_hig
+ 6.655000000e-07 V_hig
+ 6.655010000e-07 V_hig
+ 6.656000000e-07 V_hig
+ 6.656010000e-07 V_hig
+ 6.657000000e-07 V_hig
+ 6.657010000e-07 V_hig
+ 6.658000000e-07 V_hig
+ 6.658010000e-07 V_hig
+ 6.659000000e-07 V_hig
+ 6.659010000e-07 V_low
+ 6.660000000e-07 V_low
+ 6.660010000e-07 V_low
+ 6.661000000e-07 V_low
+ 6.661010000e-07 V_low
+ 6.662000000e-07 V_low
+ 6.662010000e-07 V_low
+ 6.663000000e-07 V_low
+ 6.663010000e-07 V_low
+ 6.664000000e-07 V_low
+ 6.664010000e-07 V_low
+ 6.665000000e-07 V_low
+ 6.665010000e-07 V_low
+ 6.666000000e-07 V_low
+ 6.666010000e-07 V_low
+ 6.667000000e-07 V_low
+ 6.667010000e-07 V_low
+ 6.668000000e-07 V_low
+ 6.668010000e-07 V_low
+ 6.669000000e-07 V_low
+ 6.669010000e-07 V_hig
+ 6.670000000e-07 V_hig
+ 6.670010000e-07 V_hig
+ 6.671000000e-07 V_hig
+ 6.671010000e-07 V_hig
+ 6.672000000e-07 V_hig
+ 6.672010000e-07 V_hig
+ 6.673000000e-07 V_hig
+ 6.673010000e-07 V_hig
+ 6.674000000e-07 V_hig
+ 6.674010000e-07 V_hig
+ 6.675000000e-07 V_hig
+ 6.675010000e-07 V_hig
+ 6.676000000e-07 V_hig
+ 6.676010000e-07 V_hig
+ 6.677000000e-07 V_hig
+ 6.677010000e-07 V_hig
+ 6.678000000e-07 V_hig
+ 6.678010000e-07 V_hig
+ 6.679000000e-07 V_hig
+ 6.679010000e-07 V_hig
+ 6.680000000e-07 V_hig
+ 6.680010000e-07 V_hig
+ 6.681000000e-07 V_hig
+ 6.681010000e-07 V_hig
+ 6.682000000e-07 V_hig
+ 6.682010000e-07 V_hig
+ 6.683000000e-07 V_hig
+ 6.683010000e-07 V_hig
+ 6.684000000e-07 V_hig
+ 6.684010000e-07 V_hig
+ 6.685000000e-07 V_hig
+ 6.685010000e-07 V_hig
+ 6.686000000e-07 V_hig
+ 6.686010000e-07 V_hig
+ 6.687000000e-07 V_hig
+ 6.687010000e-07 V_hig
+ 6.688000000e-07 V_hig
+ 6.688010000e-07 V_hig
+ 6.689000000e-07 V_hig
+ 6.689010000e-07 V_low
+ 6.690000000e-07 V_low
+ 6.690010000e-07 V_low
+ 6.691000000e-07 V_low
+ 6.691010000e-07 V_low
+ 6.692000000e-07 V_low
+ 6.692010000e-07 V_low
+ 6.693000000e-07 V_low
+ 6.693010000e-07 V_low
+ 6.694000000e-07 V_low
+ 6.694010000e-07 V_low
+ 6.695000000e-07 V_low
+ 6.695010000e-07 V_low
+ 6.696000000e-07 V_low
+ 6.696010000e-07 V_low
+ 6.697000000e-07 V_low
+ 6.697010000e-07 V_low
+ 6.698000000e-07 V_low
+ 6.698010000e-07 V_low
+ 6.699000000e-07 V_low
+ 6.699010000e-07 V_low
+ 6.700000000e-07 V_low
+ 6.700010000e-07 V_low
+ 6.701000000e-07 V_low
+ 6.701010000e-07 V_low
+ 6.702000000e-07 V_low
+ 6.702010000e-07 V_low
+ 6.703000000e-07 V_low
+ 6.703010000e-07 V_low
+ 6.704000000e-07 V_low
+ 6.704010000e-07 V_low
+ 6.705000000e-07 V_low
+ 6.705010000e-07 V_low
+ 6.706000000e-07 V_low
+ 6.706010000e-07 V_low
+ 6.707000000e-07 V_low
+ 6.707010000e-07 V_low
+ 6.708000000e-07 V_low
+ 6.708010000e-07 V_low
+ 6.709000000e-07 V_low
+ 6.709010000e-07 V_low
+ 6.710000000e-07 V_low
+ 6.710010000e-07 V_low
+ 6.711000000e-07 V_low
+ 6.711010000e-07 V_low
+ 6.712000000e-07 V_low
+ 6.712010000e-07 V_low
+ 6.713000000e-07 V_low
+ 6.713010000e-07 V_low
+ 6.714000000e-07 V_low
+ 6.714010000e-07 V_low
+ 6.715000000e-07 V_low
+ 6.715010000e-07 V_low
+ 6.716000000e-07 V_low
+ 6.716010000e-07 V_low
+ 6.717000000e-07 V_low
+ 6.717010000e-07 V_low
+ 6.718000000e-07 V_low
+ 6.718010000e-07 V_low
+ 6.719000000e-07 V_low
+ 6.719010000e-07 V_low
+ 6.720000000e-07 V_low
+ 6.720010000e-07 V_low
+ 6.721000000e-07 V_low
+ 6.721010000e-07 V_low
+ 6.722000000e-07 V_low
+ 6.722010000e-07 V_low
+ 6.723000000e-07 V_low
+ 6.723010000e-07 V_low
+ 6.724000000e-07 V_low
+ 6.724010000e-07 V_low
+ 6.725000000e-07 V_low
+ 6.725010000e-07 V_low
+ 6.726000000e-07 V_low
+ 6.726010000e-07 V_low
+ 6.727000000e-07 V_low
+ 6.727010000e-07 V_low
+ 6.728000000e-07 V_low
+ 6.728010000e-07 V_low
+ 6.729000000e-07 V_low
+ 6.729010000e-07 V_low
+ 6.730000000e-07 V_low
+ 6.730010000e-07 V_low
+ 6.731000000e-07 V_low
+ 6.731010000e-07 V_low
+ 6.732000000e-07 V_low
+ 6.732010000e-07 V_low
+ 6.733000000e-07 V_low
+ 6.733010000e-07 V_low
+ 6.734000000e-07 V_low
+ 6.734010000e-07 V_low
+ 6.735000000e-07 V_low
+ 6.735010000e-07 V_low
+ 6.736000000e-07 V_low
+ 6.736010000e-07 V_low
+ 6.737000000e-07 V_low
+ 6.737010000e-07 V_low
+ 6.738000000e-07 V_low
+ 6.738010000e-07 V_low
+ 6.739000000e-07 V_low
+ 6.739010000e-07 V_low
+ 6.740000000e-07 V_low
+ 6.740010000e-07 V_low
+ 6.741000000e-07 V_low
+ 6.741010000e-07 V_low
+ 6.742000000e-07 V_low
+ 6.742010000e-07 V_low
+ 6.743000000e-07 V_low
+ 6.743010000e-07 V_low
+ 6.744000000e-07 V_low
+ 6.744010000e-07 V_low
+ 6.745000000e-07 V_low
+ 6.745010000e-07 V_low
+ 6.746000000e-07 V_low
+ 6.746010000e-07 V_low
+ 6.747000000e-07 V_low
+ 6.747010000e-07 V_low
+ 6.748000000e-07 V_low
+ 6.748010000e-07 V_low
+ 6.749000000e-07 V_low
+ 6.749010000e-07 V_hig
+ 6.750000000e-07 V_hig
+ 6.750010000e-07 V_hig
+ 6.751000000e-07 V_hig
+ 6.751010000e-07 V_hig
+ 6.752000000e-07 V_hig
+ 6.752010000e-07 V_hig
+ 6.753000000e-07 V_hig
+ 6.753010000e-07 V_hig
+ 6.754000000e-07 V_hig
+ 6.754010000e-07 V_hig
+ 6.755000000e-07 V_hig
+ 6.755010000e-07 V_hig
+ 6.756000000e-07 V_hig
+ 6.756010000e-07 V_hig
+ 6.757000000e-07 V_hig
+ 6.757010000e-07 V_hig
+ 6.758000000e-07 V_hig
+ 6.758010000e-07 V_hig
+ 6.759000000e-07 V_hig
+ 6.759010000e-07 V_hig
+ 6.760000000e-07 V_hig
+ 6.760010000e-07 V_hig
+ 6.761000000e-07 V_hig
+ 6.761010000e-07 V_hig
+ 6.762000000e-07 V_hig
+ 6.762010000e-07 V_hig
+ 6.763000000e-07 V_hig
+ 6.763010000e-07 V_hig
+ 6.764000000e-07 V_hig
+ 6.764010000e-07 V_hig
+ 6.765000000e-07 V_hig
+ 6.765010000e-07 V_hig
+ 6.766000000e-07 V_hig
+ 6.766010000e-07 V_hig
+ 6.767000000e-07 V_hig
+ 6.767010000e-07 V_hig
+ 6.768000000e-07 V_hig
+ 6.768010000e-07 V_hig
+ 6.769000000e-07 V_hig
+ 6.769010000e-07 V_hig
+ 6.770000000e-07 V_hig
+ 6.770010000e-07 V_hig
+ 6.771000000e-07 V_hig
+ 6.771010000e-07 V_hig
+ 6.772000000e-07 V_hig
+ 6.772010000e-07 V_hig
+ 6.773000000e-07 V_hig
+ 6.773010000e-07 V_hig
+ 6.774000000e-07 V_hig
+ 6.774010000e-07 V_hig
+ 6.775000000e-07 V_hig
+ 6.775010000e-07 V_hig
+ 6.776000000e-07 V_hig
+ 6.776010000e-07 V_hig
+ 6.777000000e-07 V_hig
+ 6.777010000e-07 V_hig
+ 6.778000000e-07 V_hig
+ 6.778010000e-07 V_hig
+ 6.779000000e-07 V_hig
+ 6.779010000e-07 V_hig
+ 6.780000000e-07 V_hig
+ 6.780010000e-07 V_hig
+ 6.781000000e-07 V_hig
+ 6.781010000e-07 V_hig
+ 6.782000000e-07 V_hig
+ 6.782010000e-07 V_hig
+ 6.783000000e-07 V_hig
+ 6.783010000e-07 V_hig
+ 6.784000000e-07 V_hig
+ 6.784010000e-07 V_hig
+ 6.785000000e-07 V_hig
+ 6.785010000e-07 V_hig
+ 6.786000000e-07 V_hig
+ 6.786010000e-07 V_hig
+ 6.787000000e-07 V_hig
+ 6.787010000e-07 V_hig
+ 6.788000000e-07 V_hig
+ 6.788010000e-07 V_hig
+ 6.789000000e-07 V_hig
+ 6.789010000e-07 V_hig
+ 6.790000000e-07 V_hig
+ 6.790010000e-07 V_hig
+ 6.791000000e-07 V_hig
+ 6.791010000e-07 V_hig
+ 6.792000000e-07 V_hig
+ 6.792010000e-07 V_hig
+ 6.793000000e-07 V_hig
+ 6.793010000e-07 V_hig
+ 6.794000000e-07 V_hig
+ 6.794010000e-07 V_hig
+ 6.795000000e-07 V_hig
+ 6.795010000e-07 V_hig
+ 6.796000000e-07 V_hig
+ 6.796010000e-07 V_hig
+ 6.797000000e-07 V_hig
+ 6.797010000e-07 V_hig
+ 6.798000000e-07 V_hig
+ 6.798010000e-07 V_hig
+ 6.799000000e-07 V_hig
+ 6.799010000e-07 V_hig
+ 6.800000000e-07 V_hig
+ 6.800010000e-07 V_hig
+ 6.801000000e-07 V_hig
+ 6.801010000e-07 V_hig
+ 6.802000000e-07 V_hig
+ 6.802010000e-07 V_hig
+ 6.803000000e-07 V_hig
+ 6.803010000e-07 V_hig
+ 6.804000000e-07 V_hig
+ 6.804010000e-07 V_hig
+ 6.805000000e-07 V_hig
+ 6.805010000e-07 V_hig
+ 6.806000000e-07 V_hig
+ 6.806010000e-07 V_hig
+ 6.807000000e-07 V_hig
+ 6.807010000e-07 V_hig
+ 6.808000000e-07 V_hig
+ 6.808010000e-07 V_hig
+ 6.809000000e-07 V_hig
+ 6.809010000e-07 V_hig
+ 6.810000000e-07 V_hig
+ 6.810010000e-07 V_hig
+ 6.811000000e-07 V_hig
+ 6.811010000e-07 V_hig
+ 6.812000000e-07 V_hig
+ 6.812010000e-07 V_hig
+ 6.813000000e-07 V_hig
+ 6.813010000e-07 V_hig
+ 6.814000000e-07 V_hig
+ 6.814010000e-07 V_hig
+ 6.815000000e-07 V_hig
+ 6.815010000e-07 V_hig
+ 6.816000000e-07 V_hig
+ 6.816010000e-07 V_hig
+ 6.817000000e-07 V_hig
+ 6.817010000e-07 V_hig
+ 6.818000000e-07 V_hig
+ 6.818010000e-07 V_hig
+ 6.819000000e-07 V_hig
+ 6.819010000e-07 V_hig
+ 6.820000000e-07 V_hig
+ 6.820010000e-07 V_hig
+ 6.821000000e-07 V_hig
+ 6.821010000e-07 V_hig
+ 6.822000000e-07 V_hig
+ 6.822010000e-07 V_hig
+ 6.823000000e-07 V_hig
+ 6.823010000e-07 V_hig
+ 6.824000000e-07 V_hig
+ 6.824010000e-07 V_hig
+ 6.825000000e-07 V_hig
+ 6.825010000e-07 V_hig
+ 6.826000000e-07 V_hig
+ 6.826010000e-07 V_hig
+ 6.827000000e-07 V_hig
+ 6.827010000e-07 V_hig
+ 6.828000000e-07 V_hig
+ 6.828010000e-07 V_hig
+ 6.829000000e-07 V_hig
+ 6.829010000e-07 V_hig
+ 6.830000000e-07 V_hig
+ 6.830010000e-07 V_hig
+ 6.831000000e-07 V_hig
+ 6.831010000e-07 V_hig
+ 6.832000000e-07 V_hig
+ 6.832010000e-07 V_hig
+ 6.833000000e-07 V_hig
+ 6.833010000e-07 V_hig
+ 6.834000000e-07 V_hig
+ 6.834010000e-07 V_hig
+ 6.835000000e-07 V_hig
+ 6.835010000e-07 V_hig
+ 6.836000000e-07 V_hig
+ 6.836010000e-07 V_hig
+ 6.837000000e-07 V_hig
+ 6.837010000e-07 V_hig
+ 6.838000000e-07 V_hig
+ 6.838010000e-07 V_hig
+ 6.839000000e-07 V_hig
+ 6.839010000e-07 V_low
+ 6.840000000e-07 V_low
+ 6.840010000e-07 V_low
+ 6.841000000e-07 V_low
+ 6.841010000e-07 V_low
+ 6.842000000e-07 V_low
+ 6.842010000e-07 V_low
+ 6.843000000e-07 V_low
+ 6.843010000e-07 V_low
+ 6.844000000e-07 V_low
+ 6.844010000e-07 V_low
+ 6.845000000e-07 V_low
+ 6.845010000e-07 V_low
+ 6.846000000e-07 V_low
+ 6.846010000e-07 V_low
+ 6.847000000e-07 V_low
+ 6.847010000e-07 V_low
+ 6.848000000e-07 V_low
+ 6.848010000e-07 V_low
+ 6.849000000e-07 V_low
+ 6.849010000e-07 V_low
+ 6.850000000e-07 V_low
+ 6.850010000e-07 V_low
+ 6.851000000e-07 V_low
+ 6.851010000e-07 V_low
+ 6.852000000e-07 V_low
+ 6.852010000e-07 V_low
+ 6.853000000e-07 V_low
+ 6.853010000e-07 V_low
+ 6.854000000e-07 V_low
+ 6.854010000e-07 V_low
+ 6.855000000e-07 V_low
+ 6.855010000e-07 V_low
+ 6.856000000e-07 V_low
+ 6.856010000e-07 V_low
+ 6.857000000e-07 V_low
+ 6.857010000e-07 V_low
+ 6.858000000e-07 V_low
+ 6.858010000e-07 V_low
+ 6.859000000e-07 V_low
+ 6.859010000e-07 V_hig
+ 6.860000000e-07 V_hig
+ 6.860010000e-07 V_hig
+ 6.861000000e-07 V_hig
+ 6.861010000e-07 V_hig
+ 6.862000000e-07 V_hig
+ 6.862010000e-07 V_hig
+ 6.863000000e-07 V_hig
+ 6.863010000e-07 V_hig
+ 6.864000000e-07 V_hig
+ 6.864010000e-07 V_hig
+ 6.865000000e-07 V_hig
+ 6.865010000e-07 V_hig
+ 6.866000000e-07 V_hig
+ 6.866010000e-07 V_hig
+ 6.867000000e-07 V_hig
+ 6.867010000e-07 V_hig
+ 6.868000000e-07 V_hig
+ 6.868010000e-07 V_hig
+ 6.869000000e-07 V_hig
+ 6.869010000e-07 V_hig
+ 6.870000000e-07 V_hig
+ 6.870010000e-07 V_hig
+ 6.871000000e-07 V_hig
+ 6.871010000e-07 V_hig
+ 6.872000000e-07 V_hig
+ 6.872010000e-07 V_hig
+ 6.873000000e-07 V_hig
+ 6.873010000e-07 V_hig
+ 6.874000000e-07 V_hig
+ 6.874010000e-07 V_hig
+ 6.875000000e-07 V_hig
+ 6.875010000e-07 V_hig
+ 6.876000000e-07 V_hig
+ 6.876010000e-07 V_hig
+ 6.877000000e-07 V_hig
+ 6.877010000e-07 V_hig
+ 6.878000000e-07 V_hig
+ 6.878010000e-07 V_hig
+ 6.879000000e-07 V_hig
+ 6.879010000e-07 V_low
+ 6.880000000e-07 V_low
+ 6.880010000e-07 V_low
+ 6.881000000e-07 V_low
+ 6.881010000e-07 V_low
+ 6.882000000e-07 V_low
+ 6.882010000e-07 V_low
+ 6.883000000e-07 V_low
+ 6.883010000e-07 V_low
+ 6.884000000e-07 V_low
+ 6.884010000e-07 V_low
+ 6.885000000e-07 V_low
+ 6.885010000e-07 V_low
+ 6.886000000e-07 V_low
+ 6.886010000e-07 V_low
+ 6.887000000e-07 V_low
+ 6.887010000e-07 V_low
+ 6.888000000e-07 V_low
+ 6.888010000e-07 V_low
+ 6.889000000e-07 V_low
+ 6.889010000e-07 V_low
+ 6.890000000e-07 V_low
+ 6.890010000e-07 V_low
+ 6.891000000e-07 V_low
+ 6.891010000e-07 V_low
+ 6.892000000e-07 V_low
+ 6.892010000e-07 V_low
+ 6.893000000e-07 V_low
+ 6.893010000e-07 V_low
+ 6.894000000e-07 V_low
+ 6.894010000e-07 V_low
+ 6.895000000e-07 V_low
+ 6.895010000e-07 V_low
+ 6.896000000e-07 V_low
+ 6.896010000e-07 V_low
+ 6.897000000e-07 V_low
+ 6.897010000e-07 V_low
+ 6.898000000e-07 V_low
+ 6.898010000e-07 V_low
+ 6.899000000e-07 V_low
+ 6.899010000e-07 V_low
+ 6.900000000e-07 V_low
+ 6.900010000e-07 V_low
+ 6.901000000e-07 V_low
+ 6.901010000e-07 V_low
+ 6.902000000e-07 V_low
+ 6.902010000e-07 V_low
+ 6.903000000e-07 V_low
+ 6.903010000e-07 V_low
+ 6.904000000e-07 V_low
+ 6.904010000e-07 V_low
+ 6.905000000e-07 V_low
+ 6.905010000e-07 V_low
+ 6.906000000e-07 V_low
+ 6.906010000e-07 V_low
+ 6.907000000e-07 V_low
+ 6.907010000e-07 V_low
+ 6.908000000e-07 V_low
+ 6.908010000e-07 V_low
+ 6.909000000e-07 V_low
+ 6.909010000e-07 V_low
+ 6.910000000e-07 V_low
+ 6.910010000e-07 V_low
+ 6.911000000e-07 V_low
+ 6.911010000e-07 V_low
+ 6.912000000e-07 V_low
+ 6.912010000e-07 V_low
+ 6.913000000e-07 V_low
+ 6.913010000e-07 V_low
+ 6.914000000e-07 V_low
+ 6.914010000e-07 V_low
+ 6.915000000e-07 V_low
+ 6.915010000e-07 V_low
+ 6.916000000e-07 V_low
+ 6.916010000e-07 V_low
+ 6.917000000e-07 V_low
+ 6.917010000e-07 V_low
+ 6.918000000e-07 V_low
+ 6.918010000e-07 V_low
+ 6.919000000e-07 V_low
+ 6.919010000e-07 V_hig
+ 6.920000000e-07 V_hig
+ 6.920010000e-07 V_hig
+ 6.921000000e-07 V_hig
+ 6.921010000e-07 V_hig
+ 6.922000000e-07 V_hig
+ 6.922010000e-07 V_hig
+ 6.923000000e-07 V_hig
+ 6.923010000e-07 V_hig
+ 6.924000000e-07 V_hig
+ 6.924010000e-07 V_hig
+ 6.925000000e-07 V_hig
+ 6.925010000e-07 V_hig
+ 6.926000000e-07 V_hig
+ 6.926010000e-07 V_hig
+ 6.927000000e-07 V_hig
+ 6.927010000e-07 V_hig
+ 6.928000000e-07 V_hig
+ 6.928010000e-07 V_hig
+ 6.929000000e-07 V_hig
+ 6.929010000e-07 V_hig
+ 6.930000000e-07 V_hig
+ 6.930010000e-07 V_hig
+ 6.931000000e-07 V_hig
+ 6.931010000e-07 V_hig
+ 6.932000000e-07 V_hig
+ 6.932010000e-07 V_hig
+ 6.933000000e-07 V_hig
+ 6.933010000e-07 V_hig
+ 6.934000000e-07 V_hig
+ 6.934010000e-07 V_hig
+ 6.935000000e-07 V_hig
+ 6.935010000e-07 V_hig
+ 6.936000000e-07 V_hig
+ 6.936010000e-07 V_hig
+ 6.937000000e-07 V_hig
+ 6.937010000e-07 V_hig
+ 6.938000000e-07 V_hig
+ 6.938010000e-07 V_hig
+ 6.939000000e-07 V_hig
+ 6.939010000e-07 V_hig
+ 6.940000000e-07 V_hig
+ 6.940010000e-07 V_hig
+ 6.941000000e-07 V_hig
+ 6.941010000e-07 V_hig
+ 6.942000000e-07 V_hig
+ 6.942010000e-07 V_hig
+ 6.943000000e-07 V_hig
+ 6.943010000e-07 V_hig
+ 6.944000000e-07 V_hig
+ 6.944010000e-07 V_hig
+ 6.945000000e-07 V_hig
+ 6.945010000e-07 V_hig
+ 6.946000000e-07 V_hig
+ 6.946010000e-07 V_hig
+ 6.947000000e-07 V_hig
+ 6.947010000e-07 V_hig
+ 6.948000000e-07 V_hig
+ 6.948010000e-07 V_hig
+ 6.949000000e-07 V_hig
+ 6.949010000e-07 V_low
+ 6.950000000e-07 V_low
+ 6.950010000e-07 V_low
+ 6.951000000e-07 V_low
+ 6.951010000e-07 V_low
+ 6.952000000e-07 V_low
+ 6.952010000e-07 V_low
+ 6.953000000e-07 V_low
+ 6.953010000e-07 V_low
+ 6.954000000e-07 V_low
+ 6.954010000e-07 V_low
+ 6.955000000e-07 V_low
+ 6.955010000e-07 V_low
+ 6.956000000e-07 V_low
+ 6.956010000e-07 V_low
+ 6.957000000e-07 V_low
+ 6.957010000e-07 V_low
+ 6.958000000e-07 V_low
+ 6.958010000e-07 V_low
+ 6.959000000e-07 V_low
+ 6.959010000e-07 V_low
+ 6.960000000e-07 V_low
+ 6.960010000e-07 V_low
+ 6.961000000e-07 V_low
+ 6.961010000e-07 V_low
+ 6.962000000e-07 V_low
+ 6.962010000e-07 V_low
+ 6.963000000e-07 V_low
+ 6.963010000e-07 V_low
+ 6.964000000e-07 V_low
+ 6.964010000e-07 V_low
+ 6.965000000e-07 V_low
+ 6.965010000e-07 V_low
+ 6.966000000e-07 V_low
+ 6.966010000e-07 V_low
+ 6.967000000e-07 V_low
+ 6.967010000e-07 V_low
+ 6.968000000e-07 V_low
+ 6.968010000e-07 V_low
+ 6.969000000e-07 V_low
+ 6.969010000e-07 V_hig
+ 6.970000000e-07 V_hig
+ 6.970010000e-07 V_hig
+ 6.971000000e-07 V_hig
+ 6.971010000e-07 V_hig
+ 6.972000000e-07 V_hig
+ 6.972010000e-07 V_hig
+ 6.973000000e-07 V_hig
+ 6.973010000e-07 V_hig
+ 6.974000000e-07 V_hig
+ 6.974010000e-07 V_hig
+ 6.975000000e-07 V_hig
+ 6.975010000e-07 V_hig
+ 6.976000000e-07 V_hig
+ 6.976010000e-07 V_hig
+ 6.977000000e-07 V_hig
+ 6.977010000e-07 V_hig
+ 6.978000000e-07 V_hig
+ 6.978010000e-07 V_hig
+ 6.979000000e-07 V_hig
+ 6.979010000e-07 V_hig
+ 6.980000000e-07 V_hig
+ 6.980010000e-07 V_hig
+ 6.981000000e-07 V_hig
+ 6.981010000e-07 V_hig
+ 6.982000000e-07 V_hig
+ 6.982010000e-07 V_hig
+ 6.983000000e-07 V_hig
+ 6.983010000e-07 V_hig
+ 6.984000000e-07 V_hig
+ 6.984010000e-07 V_hig
+ 6.985000000e-07 V_hig
+ 6.985010000e-07 V_hig
+ 6.986000000e-07 V_hig
+ 6.986010000e-07 V_hig
+ 6.987000000e-07 V_hig
+ 6.987010000e-07 V_hig
+ 6.988000000e-07 V_hig
+ 6.988010000e-07 V_hig
+ 6.989000000e-07 V_hig
+ 6.989010000e-07 V_hig
+ 6.990000000e-07 V_hig
+ 6.990010000e-07 V_hig
+ 6.991000000e-07 V_hig
+ 6.991010000e-07 V_hig
+ 6.992000000e-07 V_hig
+ 6.992010000e-07 V_hig
+ 6.993000000e-07 V_hig
+ 6.993010000e-07 V_hig
+ 6.994000000e-07 V_hig
+ 6.994010000e-07 V_hig
+ 6.995000000e-07 V_hig
+ 6.995010000e-07 V_hig
+ 6.996000000e-07 V_hig
+ 6.996010000e-07 V_hig
+ 6.997000000e-07 V_hig
+ 6.997010000e-07 V_hig
+ 6.998000000e-07 V_hig
+ 6.998010000e-07 V_hig
+ 6.999000000e-07 V_hig
+ 6.999010000e-07 V_low
+ 7.000000000e-07 V_low
+ 7.000010000e-07 V_low
+ 7.001000000e-07 V_low
+ 7.001010000e-07 V_low
+ 7.002000000e-07 V_low
+ 7.002010000e-07 V_low
+ 7.003000000e-07 V_low
+ 7.003010000e-07 V_low
+ 7.004000000e-07 V_low
+ 7.004010000e-07 V_low
+ 7.005000000e-07 V_low
+ 7.005010000e-07 V_low
+ 7.006000000e-07 V_low
+ 7.006010000e-07 V_low
+ 7.007000000e-07 V_low
+ 7.007010000e-07 V_low
+ 7.008000000e-07 V_low
+ 7.008010000e-07 V_low
+ 7.009000000e-07 V_low
+ 7.009010000e-07 V_low
+ 7.010000000e-07 V_low
+ 7.010010000e-07 V_low
+ 7.011000000e-07 V_low
+ 7.011010000e-07 V_low
+ 7.012000000e-07 V_low
+ 7.012010000e-07 V_low
+ 7.013000000e-07 V_low
+ 7.013010000e-07 V_low
+ 7.014000000e-07 V_low
+ 7.014010000e-07 V_low
+ 7.015000000e-07 V_low
+ 7.015010000e-07 V_low
+ 7.016000000e-07 V_low
+ 7.016010000e-07 V_low
+ 7.017000000e-07 V_low
+ 7.017010000e-07 V_low
+ 7.018000000e-07 V_low
+ 7.018010000e-07 V_low
+ 7.019000000e-07 V_low
+ 7.019010000e-07 V_hig
+ 7.020000000e-07 V_hig
+ 7.020010000e-07 V_hig
+ 7.021000000e-07 V_hig
+ 7.021010000e-07 V_hig
+ 7.022000000e-07 V_hig
+ 7.022010000e-07 V_hig
+ 7.023000000e-07 V_hig
+ 7.023010000e-07 V_hig
+ 7.024000000e-07 V_hig
+ 7.024010000e-07 V_hig
+ 7.025000000e-07 V_hig
+ 7.025010000e-07 V_hig
+ 7.026000000e-07 V_hig
+ 7.026010000e-07 V_hig
+ 7.027000000e-07 V_hig
+ 7.027010000e-07 V_hig
+ 7.028000000e-07 V_hig
+ 7.028010000e-07 V_hig
+ 7.029000000e-07 V_hig
+ 7.029010000e-07 V_hig
+ 7.030000000e-07 V_hig
+ 7.030010000e-07 V_hig
+ 7.031000000e-07 V_hig
+ 7.031010000e-07 V_hig
+ 7.032000000e-07 V_hig
+ 7.032010000e-07 V_hig
+ 7.033000000e-07 V_hig
+ 7.033010000e-07 V_hig
+ 7.034000000e-07 V_hig
+ 7.034010000e-07 V_hig
+ 7.035000000e-07 V_hig
+ 7.035010000e-07 V_hig
+ 7.036000000e-07 V_hig
+ 7.036010000e-07 V_hig
+ 7.037000000e-07 V_hig
+ 7.037010000e-07 V_hig
+ 7.038000000e-07 V_hig
+ 7.038010000e-07 V_hig
+ 7.039000000e-07 V_hig
+ 7.039010000e-07 V_hig
+ 7.040000000e-07 V_hig
+ 7.040010000e-07 V_hig
+ 7.041000000e-07 V_hig
+ 7.041010000e-07 V_hig
+ 7.042000000e-07 V_hig
+ 7.042010000e-07 V_hig
+ 7.043000000e-07 V_hig
+ 7.043010000e-07 V_hig
+ 7.044000000e-07 V_hig
+ 7.044010000e-07 V_hig
+ 7.045000000e-07 V_hig
+ 7.045010000e-07 V_hig
+ 7.046000000e-07 V_hig
+ 7.046010000e-07 V_hig
+ 7.047000000e-07 V_hig
+ 7.047010000e-07 V_hig
+ 7.048000000e-07 V_hig
+ 7.048010000e-07 V_hig
+ 7.049000000e-07 V_hig
+ 7.049010000e-07 V_low
+ 7.050000000e-07 V_low
+ 7.050010000e-07 V_low
+ 7.051000000e-07 V_low
+ 7.051010000e-07 V_low
+ 7.052000000e-07 V_low
+ 7.052010000e-07 V_low
+ 7.053000000e-07 V_low
+ 7.053010000e-07 V_low
+ 7.054000000e-07 V_low
+ 7.054010000e-07 V_low
+ 7.055000000e-07 V_low
+ 7.055010000e-07 V_low
+ 7.056000000e-07 V_low
+ 7.056010000e-07 V_low
+ 7.057000000e-07 V_low
+ 7.057010000e-07 V_low
+ 7.058000000e-07 V_low
+ 7.058010000e-07 V_low
+ 7.059000000e-07 V_low
+ 7.059010000e-07 V_low
+ 7.060000000e-07 V_low
+ 7.060010000e-07 V_low
+ 7.061000000e-07 V_low
+ 7.061010000e-07 V_low
+ 7.062000000e-07 V_low
+ 7.062010000e-07 V_low
+ 7.063000000e-07 V_low
+ 7.063010000e-07 V_low
+ 7.064000000e-07 V_low
+ 7.064010000e-07 V_low
+ 7.065000000e-07 V_low
+ 7.065010000e-07 V_low
+ 7.066000000e-07 V_low
+ 7.066010000e-07 V_low
+ 7.067000000e-07 V_low
+ 7.067010000e-07 V_low
+ 7.068000000e-07 V_low
+ 7.068010000e-07 V_low
+ 7.069000000e-07 V_low
+ 7.069010000e-07 V_hig
+ 7.070000000e-07 V_hig
+ 7.070010000e-07 V_hig
+ 7.071000000e-07 V_hig
+ 7.071010000e-07 V_hig
+ 7.072000000e-07 V_hig
+ 7.072010000e-07 V_hig
+ 7.073000000e-07 V_hig
+ 7.073010000e-07 V_hig
+ 7.074000000e-07 V_hig
+ 7.074010000e-07 V_hig
+ 7.075000000e-07 V_hig
+ 7.075010000e-07 V_hig
+ 7.076000000e-07 V_hig
+ 7.076010000e-07 V_hig
+ 7.077000000e-07 V_hig
+ 7.077010000e-07 V_hig
+ 7.078000000e-07 V_hig
+ 7.078010000e-07 V_hig
+ 7.079000000e-07 V_hig
+ 7.079010000e-07 V_low
+ 7.080000000e-07 V_low
+ 7.080010000e-07 V_low
+ 7.081000000e-07 V_low
+ 7.081010000e-07 V_low
+ 7.082000000e-07 V_low
+ 7.082010000e-07 V_low
+ 7.083000000e-07 V_low
+ 7.083010000e-07 V_low
+ 7.084000000e-07 V_low
+ 7.084010000e-07 V_low
+ 7.085000000e-07 V_low
+ 7.085010000e-07 V_low
+ 7.086000000e-07 V_low
+ 7.086010000e-07 V_low
+ 7.087000000e-07 V_low
+ 7.087010000e-07 V_low
+ 7.088000000e-07 V_low
+ 7.088010000e-07 V_low
+ 7.089000000e-07 V_low
+ 7.089010000e-07 V_low
+ 7.090000000e-07 V_low
+ 7.090010000e-07 V_low
+ 7.091000000e-07 V_low
+ 7.091010000e-07 V_low
+ 7.092000000e-07 V_low
+ 7.092010000e-07 V_low
+ 7.093000000e-07 V_low
+ 7.093010000e-07 V_low
+ 7.094000000e-07 V_low
+ 7.094010000e-07 V_low
+ 7.095000000e-07 V_low
+ 7.095010000e-07 V_low
+ 7.096000000e-07 V_low
+ 7.096010000e-07 V_low
+ 7.097000000e-07 V_low
+ 7.097010000e-07 V_low
+ 7.098000000e-07 V_low
+ 7.098010000e-07 V_low
+ 7.099000000e-07 V_low
+ 7.099010000e-07 V_hig
+ 7.100000000e-07 V_hig
+ 7.100010000e-07 V_hig
+ 7.101000000e-07 V_hig
+ 7.101010000e-07 V_hig
+ 7.102000000e-07 V_hig
+ 7.102010000e-07 V_hig
+ 7.103000000e-07 V_hig
+ 7.103010000e-07 V_hig
+ 7.104000000e-07 V_hig
+ 7.104010000e-07 V_hig
+ 7.105000000e-07 V_hig
+ 7.105010000e-07 V_hig
+ 7.106000000e-07 V_hig
+ 7.106010000e-07 V_hig
+ 7.107000000e-07 V_hig
+ 7.107010000e-07 V_hig
+ 7.108000000e-07 V_hig
+ 7.108010000e-07 V_hig
+ 7.109000000e-07 V_hig
+ 7.109010000e-07 V_hig
+ 7.110000000e-07 V_hig
+ 7.110010000e-07 V_hig
+ 7.111000000e-07 V_hig
+ 7.111010000e-07 V_hig
+ 7.112000000e-07 V_hig
+ 7.112010000e-07 V_hig
+ 7.113000000e-07 V_hig
+ 7.113010000e-07 V_hig
+ 7.114000000e-07 V_hig
+ 7.114010000e-07 V_hig
+ 7.115000000e-07 V_hig
+ 7.115010000e-07 V_hig
+ 7.116000000e-07 V_hig
+ 7.116010000e-07 V_hig
+ 7.117000000e-07 V_hig
+ 7.117010000e-07 V_hig
+ 7.118000000e-07 V_hig
+ 7.118010000e-07 V_hig
+ 7.119000000e-07 V_hig
+ 7.119010000e-07 V_low
+ 7.120000000e-07 V_low
+ 7.120010000e-07 V_low
+ 7.121000000e-07 V_low
+ 7.121010000e-07 V_low
+ 7.122000000e-07 V_low
+ 7.122010000e-07 V_low
+ 7.123000000e-07 V_low
+ 7.123010000e-07 V_low
+ 7.124000000e-07 V_low
+ 7.124010000e-07 V_low
+ 7.125000000e-07 V_low
+ 7.125010000e-07 V_low
+ 7.126000000e-07 V_low
+ 7.126010000e-07 V_low
+ 7.127000000e-07 V_low
+ 7.127010000e-07 V_low
+ 7.128000000e-07 V_low
+ 7.128010000e-07 V_low
+ 7.129000000e-07 V_low
+ 7.129010000e-07 V_hig
+ 7.130000000e-07 V_hig
+ 7.130010000e-07 V_hig
+ 7.131000000e-07 V_hig
+ 7.131010000e-07 V_hig
+ 7.132000000e-07 V_hig
+ 7.132010000e-07 V_hig
+ 7.133000000e-07 V_hig
+ 7.133010000e-07 V_hig
+ 7.134000000e-07 V_hig
+ 7.134010000e-07 V_hig
+ 7.135000000e-07 V_hig
+ 7.135010000e-07 V_hig
+ 7.136000000e-07 V_hig
+ 7.136010000e-07 V_hig
+ 7.137000000e-07 V_hig
+ 7.137010000e-07 V_hig
+ 7.138000000e-07 V_hig
+ 7.138010000e-07 V_hig
+ 7.139000000e-07 V_hig
+ 7.139010000e-07 V_low
+ 7.140000000e-07 V_low
+ 7.140010000e-07 V_low
+ 7.141000000e-07 V_low
+ 7.141010000e-07 V_low
+ 7.142000000e-07 V_low
+ 7.142010000e-07 V_low
+ 7.143000000e-07 V_low
+ 7.143010000e-07 V_low
+ 7.144000000e-07 V_low
+ 7.144010000e-07 V_low
+ 7.145000000e-07 V_low
+ 7.145010000e-07 V_low
+ 7.146000000e-07 V_low
+ 7.146010000e-07 V_low
+ 7.147000000e-07 V_low
+ 7.147010000e-07 V_low
+ 7.148000000e-07 V_low
+ 7.148010000e-07 V_low
+ 7.149000000e-07 V_low
+ 7.149010000e-07 V_hig
+ 7.150000000e-07 V_hig
+ 7.150010000e-07 V_hig
+ 7.151000000e-07 V_hig
+ 7.151010000e-07 V_hig
+ 7.152000000e-07 V_hig
+ 7.152010000e-07 V_hig
+ 7.153000000e-07 V_hig
+ 7.153010000e-07 V_hig
+ 7.154000000e-07 V_hig
+ 7.154010000e-07 V_hig
+ 7.155000000e-07 V_hig
+ 7.155010000e-07 V_hig
+ 7.156000000e-07 V_hig
+ 7.156010000e-07 V_hig
+ 7.157000000e-07 V_hig
+ 7.157010000e-07 V_hig
+ 7.158000000e-07 V_hig
+ 7.158010000e-07 V_hig
+ 7.159000000e-07 V_hig
+ 7.159010000e-07 V_hig
+ 7.160000000e-07 V_hig
+ 7.160010000e-07 V_hig
+ 7.161000000e-07 V_hig
+ 7.161010000e-07 V_hig
+ 7.162000000e-07 V_hig
+ 7.162010000e-07 V_hig
+ 7.163000000e-07 V_hig
+ 7.163010000e-07 V_hig
+ 7.164000000e-07 V_hig
+ 7.164010000e-07 V_hig
+ 7.165000000e-07 V_hig
+ 7.165010000e-07 V_hig
+ 7.166000000e-07 V_hig
+ 7.166010000e-07 V_hig
+ 7.167000000e-07 V_hig
+ 7.167010000e-07 V_hig
+ 7.168000000e-07 V_hig
+ 7.168010000e-07 V_hig
+ 7.169000000e-07 V_hig
+ 7.169010000e-07 V_hig
+ 7.170000000e-07 V_hig
+ 7.170010000e-07 V_hig
+ 7.171000000e-07 V_hig
+ 7.171010000e-07 V_hig
+ 7.172000000e-07 V_hig
+ 7.172010000e-07 V_hig
+ 7.173000000e-07 V_hig
+ 7.173010000e-07 V_hig
+ 7.174000000e-07 V_hig
+ 7.174010000e-07 V_hig
+ 7.175000000e-07 V_hig
+ 7.175010000e-07 V_hig
+ 7.176000000e-07 V_hig
+ 7.176010000e-07 V_hig
+ 7.177000000e-07 V_hig
+ 7.177010000e-07 V_hig
+ 7.178000000e-07 V_hig
+ 7.178010000e-07 V_hig
+ 7.179000000e-07 V_hig
+ 7.179010000e-07 V_low
+ 7.180000000e-07 V_low
+ 7.180010000e-07 V_low
+ 7.181000000e-07 V_low
+ 7.181010000e-07 V_low
+ 7.182000000e-07 V_low
+ 7.182010000e-07 V_low
+ 7.183000000e-07 V_low
+ 7.183010000e-07 V_low
+ 7.184000000e-07 V_low
+ 7.184010000e-07 V_low
+ 7.185000000e-07 V_low
+ 7.185010000e-07 V_low
+ 7.186000000e-07 V_low
+ 7.186010000e-07 V_low
+ 7.187000000e-07 V_low
+ 7.187010000e-07 V_low
+ 7.188000000e-07 V_low
+ 7.188010000e-07 V_low
+ 7.189000000e-07 V_low
+ 7.189010000e-07 V_low
+ 7.190000000e-07 V_low
+ 7.190010000e-07 V_low
+ 7.191000000e-07 V_low
+ 7.191010000e-07 V_low
+ 7.192000000e-07 V_low
+ 7.192010000e-07 V_low
+ 7.193000000e-07 V_low
+ 7.193010000e-07 V_low
+ 7.194000000e-07 V_low
+ 7.194010000e-07 V_low
+ 7.195000000e-07 V_low
+ 7.195010000e-07 V_low
+ 7.196000000e-07 V_low
+ 7.196010000e-07 V_low
+ 7.197000000e-07 V_low
+ 7.197010000e-07 V_low
+ 7.198000000e-07 V_low
+ 7.198010000e-07 V_low
+ 7.199000000e-07 V_low
+ 7.199010000e-07 V_low
+ 7.200000000e-07 V_low
+ 7.200010000e-07 V_low
+ 7.201000000e-07 V_low
+ 7.201010000e-07 V_low
+ 7.202000000e-07 V_low
+ 7.202010000e-07 V_low
+ 7.203000000e-07 V_low
+ 7.203010000e-07 V_low
+ 7.204000000e-07 V_low
+ 7.204010000e-07 V_low
+ 7.205000000e-07 V_low
+ 7.205010000e-07 V_low
+ 7.206000000e-07 V_low
+ 7.206010000e-07 V_low
+ 7.207000000e-07 V_low
+ 7.207010000e-07 V_low
+ 7.208000000e-07 V_low
+ 7.208010000e-07 V_low
+ 7.209000000e-07 V_low
+ 7.209010000e-07 V_low
+ 7.210000000e-07 V_low
+ 7.210010000e-07 V_low
+ 7.211000000e-07 V_low
+ 7.211010000e-07 V_low
+ 7.212000000e-07 V_low
+ 7.212010000e-07 V_low
+ 7.213000000e-07 V_low
+ 7.213010000e-07 V_low
+ 7.214000000e-07 V_low
+ 7.214010000e-07 V_low
+ 7.215000000e-07 V_low
+ 7.215010000e-07 V_low
+ 7.216000000e-07 V_low
+ 7.216010000e-07 V_low
+ 7.217000000e-07 V_low
+ 7.217010000e-07 V_low
+ 7.218000000e-07 V_low
+ 7.218010000e-07 V_low
+ 7.219000000e-07 V_low
+ 7.219010000e-07 V_hig
+ 7.220000000e-07 V_hig
+ 7.220010000e-07 V_hig
+ 7.221000000e-07 V_hig
+ 7.221010000e-07 V_hig
+ 7.222000000e-07 V_hig
+ 7.222010000e-07 V_hig
+ 7.223000000e-07 V_hig
+ 7.223010000e-07 V_hig
+ 7.224000000e-07 V_hig
+ 7.224010000e-07 V_hig
+ 7.225000000e-07 V_hig
+ 7.225010000e-07 V_hig
+ 7.226000000e-07 V_hig
+ 7.226010000e-07 V_hig
+ 7.227000000e-07 V_hig
+ 7.227010000e-07 V_hig
+ 7.228000000e-07 V_hig
+ 7.228010000e-07 V_hig
+ 7.229000000e-07 V_hig
+ 7.229010000e-07 V_hig
+ 7.230000000e-07 V_hig
+ 7.230010000e-07 V_hig
+ 7.231000000e-07 V_hig
+ 7.231010000e-07 V_hig
+ 7.232000000e-07 V_hig
+ 7.232010000e-07 V_hig
+ 7.233000000e-07 V_hig
+ 7.233010000e-07 V_hig
+ 7.234000000e-07 V_hig
+ 7.234010000e-07 V_hig
+ 7.235000000e-07 V_hig
+ 7.235010000e-07 V_hig
+ 7.236000000e-07 V_hig
+ 7.236010000e-07 V_hig
+ 7.237000000e-07 V_hig
+ 7.237010000e-07 V_hig
+ 7.238000000e-07 V_hig
+ 7.238010000e-07 V_hig
+ 7.239000000e-07 V_hig
+ 7.239010000e-07 V_hig
+ 7.240000000e-07 V_hig
+ 7.240010000e-07 V_hig
+ 7.241000000e-07 V_hig
+ 7.241010000e-07 V_hig
+ 7.242000000e-07 V_hig
+ 7.242010000e-07 V_hig
+ 7.243000000e-07 V_hig
+ 7.243010000e-07 V_hig
+ 7.244000000e-07 V_hig
+ 7.244010000e-07 V_hig
+ 7.245000000e-07 V_hig
+ 7.245010000e-07 V_hig
+ 7.246000000e-07 V_hig
+ 7.246010000e-07 V_hig
+ 7.247000000e-07 V_hig
+ 7.247010000e-07 V_hig
+ 7.248000000e-07 V_hig
+ 7.248010000e-07 V_hig
+ 7.249000000e-07 V_hig
+ 7.249010000e-07 V_hig
+ 7.250000000e-07 V_hig
+ 7.250010000e-07 V_hig
+ 7.251000000e-07 V_hig
+ 7.251010000e-07 V_hig
+ 7.252000000e-07 V_hig
+ 7.252010000e-07 V_hig
+ 7.253000000e-07 V_hig
+ 7.253010000e-07 V_hig
+ 7.254000000e-07 V_hig
+ 7.254010000e-07 V_hig
+ 7.255000000e-07 V_hig
+ 7.255010000e-07 V_hig
+ 7.256000000e-07 V_hig
+ 7.256010000e-07 V_hig
+ 7.257000000e-07 V_hig
+ 7.257010000e-07 V_hig
+ 7.258000000e-07 V_hig
+ 7.258010000e-07 V_hig
+ 7.259000000e-07 V_hig
+ 7.259010000e-07 V_low
+ 7.260000000e-07 V_low
+ 7.260010000e-07 V_low
+ 7.261000000e-07 V_low
+ 7.261010000e-07 V_low
+ 7.262000000e-07 V_low
+ 7.262010000e-07 V_low
+ 7.263000000e-07 V_low
+ 7.263010000e-07 V_low
+ 7.264000000e-07 V_low
+ 7.264010000e-07 V_low
+ 7.265000000e-07 V_low
+ 7.265010000e-07 V_low
+ 7.266000000e-07 V_low
+ 7.266010000e-07 V_low
+ 7.267000000e-07 V_low
+ 7.267010000e-07 V_low
+ 7.268000000e-07 V_low
+ 7.268010000e-07 V_low
+ 7.269000000e-07 V_low
+ 7.269010000e-07 V_low
+ 7.270000000e-07 V_low
+ 7.270010000e-07 V_low
+ 7.271000000e-07 V_low
+ 7.271010000e-07 V_low
+ 7.272000000e-07 V_low
+ 7.272010000e-07 V_low
+ 7.273000000e-07 V_low
+ 7.273010000e-07 V_low
+ 7.274000000e-07 V_low
+ 7.274010000e-07 V_low
+ 7.275000000e-07 V_low
+ 7.275010000e-07 V_low
+ 7.276000000e-07 V_low
+ 7.276010000e-07 V_low
+ 7.277000000e-07 V_low
+ 7.277010000e-07 V_low
+ 7.278000000e-07 V_low
+ 7.278010000e-07 V_low
+ 7.279000000e-07 V_low
+ 7.279010000e-07 V_hig
+ 7.280000000e-07 V_hig
+ 7.280010000e-07 V_hig
+ 7.281000000e-07 V_hig
+ 7.281010000e-07 V_hig
+ 7.282000000e-07 V_hig
+ 7.282010000e-07 V_hig
+ 7.283000000e-07 V_hig
+ 7.283010000e-07 V_hig
+ 7.284000000e-07 V_hig
+ 7.284010000e-07 V_hig
+ 7.285000000e-07 V_hig
+ 7.285010000e-07 V_hig
+ 7.286000000e-07 V_hig
+ 7.286010000e-07 V_hig
+ 7.287000000e-07 V_hig
+ 7.287010000e-07 V_hig
+ 7.288000000e-07 V_hig
+ 7.288010000e-07 V_hig
+ 7.289000000e-07 V_hig
+ 7.289010000e-07 V_low
+ 7.290000000e-07 V_low
+ 7.290010000e-07 V_low
+ 7.291000000e-07 V_low
+ 7.291010000e-07 V_low
+ 7.292000000e-07 V_low
+ 7.292010000e-07 V_low
+ 7.293000000e-07 V_low
+ 7.293010000e-07 V_low
+ 7.294000000e-07 V_low
+ 7.294010000e-07 V_low
+ 7.295000000e-07 V_low
+ 7.295010000e-07 V_low
+ 7.296000000e-07 V_low
+ 7.296010000e-07 V_low
+ 7.297000000e-07 V_low
+ 7.297010000e-07 V_low
+ 7.298000000e-07 V_low
+ 7.298010000e-07 V_low
+ 7.299000000e-07 V_low
+ 7.299010000e-07 V_hig
+ 7.300000000e-07 V_hig
+ 7.300010000e-07 V_hig
+ 7.301000000e-07 V_hig
+ 7.301010000e-07 V_hig
+ 7.302000000e-07 V_hig
+ 7.302010000e-07 V_hig
+ 7.303000000e-07 V_hig
+ 7.303010000e-07 V_hig
+ 7.304000000e-07 V_hig
+ 7.304010000e-07 V_hig
+ 7.305000000e-07 V_hig
+ 7.305010000e-07 V_hig
+ 7.306000000e-07 V_hig
+ 7.306010000e-07 V_hig
+ 7.307000000e-07 V_hig
+ 7.307010000e-07 V_hig
+ 7.308000000e-07 V_hig
+ 7.308010000e-07 V_hig
+ 7.309000000e-07 V_hig
+ 7.309010000e-07 V_hig
+ 7.310000000e-07 V_hig
+ 7.310010000e-07 V_hig
+ 7.311000000e-07 V_hig
+ 7.311010000e-07 V_hig
+ 7.312000000e-07 V_hig
+ 7.312010000e-07 V_hig
+ 7.313000000e-07 V_hig
+ 7.313010000e-07 V_hig
+ 7.314000000e-07 V_hig
+ 7.314010000e-07 V_hig
+ 7.315000000e-07 V_hig
+ 7.315010000e-07 V_hig
+ 7.316000000e-07 V_hig
+ 7.316010000e-07 V_hig
+ 7.317000000e-07 V_hig
+ 7.317010000e-07 V_hig
+ 7.318000000e-07 V_hig
+ 7.318010000e-07 V_hig
+ 7.319000000e-07 V_hig
+ 7.319010000e-07 V_low
+ 7.320000000e-07 V_low
+ 7.320010000e-07 V_low
+ 7.321000000e-07 V_low
+ 7.321010000e-07 V_low
+ 7.322000000e-07 V_low
+ 7.322010000e-07 V_low
+ 7.323000000e-07 V_low
+ 7.323010000e-07 V_low
+ 7.324000000e-07 V_low
+ 7.324010000e-07 V_low
+ 7.325000000e-07 V_low
+ 7.325010000e-07 V_low
+ 7.326000000e-07 V_low
+ 7.326010000e-07 V_low
+ 7.327000000e-07 V_low
+ 7.327010000e-07 V_low
+ 7.328000000e-07 V_low
+ 7.328010000e-07 V_low
+ 7.329000000e-07 V_low
+ 7.329010000e-07 V_hig
+ 7.330000000e-07 V_hig
+ 7.330010000e-07 V_hig
+ 7.331000000e-07 V_hig
+ 7.331010000e-07 V_hig
+ 7.332000000e-07 V_hig
+ 7.332010000e-07 V_hig
+ 7.333000000e-07 V_hig
+ 7.333010000e-07 V_hig
+ 7.334000000e-07 V_hig
+ 7.334010000e-07 V_hig
+ 7.335000000e-07 V_hig
+ 7.335010000e-07 V_hig
+ 7.336000000e-07 V_hig
+ 7.336010000e-07 V_hig
+ 7.337000000e-07 V_hig
+ 7.337010000e-07 V_hig
+ 7.338000000e-07 V_hig
+ 7.338010000e-07 V_hig
+ 7.339000000e-07 V_hig
+ 7.339010000e-07 V_hig
+ 7.340000000e-07 V_hig
+ 7.340010000e-07 V_hig
+ 7.341000000e-07 V_hig
+ 7.341010000e-07 V_hig
+ 7.342000000e-07 V_hig
+ 7.342010000e-07 V_hig
+ 7.343000000e-07 V_hig
+ 7.343010000e-07 V_hig
+ 7.344000000e-07 V_hig
+ 7.344010000e-07 V_hig
+ 7.345000000e-07 V_hig
+ 7.345010000e-07 V_hig
+ 7.346000000e-07 V_hig
+ 7.346010000e-07 V_hig
+ 7.347000000e-07 V_hig
+ 7.347010000e-07 V_hig
+ 7.348000000e-07 V_hig
+ 7.348010000e-07 V_hig
+ 7.349000000e-07 V_hig
+ 7.349010000e-07 V_low
+ 7.350000000e-07 V_low
+ 7.350010000e-07 V_low
+ 7.351000000e-07 V_low
+ 7.351010000e-07 V_low
+ 7.352000000e-07 V_low
+ 7.352010000e-07 V_low
+ 7.353000000e-07 V_low
+ 7.353010000e-07 V_low
+ 7.354000000e-07 V_low
+ 7.354010000e-07 V_low
+ 7.355000000e-07 V_low
+ 7.355010000e-07 V_low
+ 7.356000000e-07 V_low
+ 7.356010000e-07 V_low
+ 7.357000000e-07 V_low
+ 7.357010000e-07 V_low
+ 7.358000000e-07 V_low
+ 7.358010000e-07 V_low
+ 7.359000000e-07 V_low
+ 7.359010000e-07 V_low
+ 7.360000000e-07 V_low
+ 7.360010000e-07 V_low
+ 7.361000000e-07 V_low
+ 7.361010000e-07 V_low
+ 7.362000000e-07 V_low
+ 7.362010000e-07 V_low
+ 7.363000000e-07 V_low
+ 7.363010000e-07 V_low
+ 7.364000000e-07 V_low
+ 7.364010000e-07 V_low
+ 7.365000000e-07 V_low
+ 7.365010000e-07 V_low
+ 7.366000000e-07 V_low
+ 7.366010000e-07 V_low
+ 7.367000000e-07 V_low
+ 7.367010000e-07 V_low
+ 7.368000000e-07 V_low
+ 7.368010000e-07 V_low
+ 7.369000000e-07 V_low
+ 7.369010000e-07 V_hig
+ 7.370000000e-07 V_hig
+ 7.370010000e-07 V_hig
+ 7.371000000e-07 V_hig
+ 7.371010000e-07 V_hig
+ 7.372000000e-07 V_hig
+ 7.372010000e-07 V_hig
+ 7.373000000e-07 V_hig
+ 7.373010000e-07 V_hig
+ 7.374000000e-07 V_hig
+ 7.374010000e-07 V_hig
+ 7.375000000e-07 V_hig
+ 7.375010000e-07 V_hig
+ 7.376000000e-07 V_hig
+ 7.376010000e-07 V_hig
+ 7.377000000e-07 V_hig
+ 7.377010000e-07 V_hig
+ 7.378000000e-07 V_hig
+ 7.378010000e-07 V_hig
+ 7.379000000e-07 V_hig
+ 7.379010000e-07 V_hig
+ 7.380000000e-07 V_hig
+ 7.380010000e-07 V_hig
+ 7.381000000e-07 V_hig
+ 7.381010000e-07 V_hig
+ 7.382000000e-07 V_hig
+ 7.382010000e-07 V_hig
+ 7.383000000e-07 V_hig
+ 7.383010000e-07 V_hig
+ 7.384000000e-07 V_hig
+ 7.384010000e-07 V_hig
+ 7.385000000e-07 V_hig
+ 7.385010000e-07 V_hig
+ 7.386000000e-07 V_hig
+ 7.386010000e-07 V_hig
+ 7.387000000e-07 V_hig
+ 7.387010000e-07 V_hig
+ 7.388000000e-07 V_hig
+ 7.388010000e-07 V_hig
+ 7.389000000e-07 V_hig
+ 7.389010000e-07 V_low
+ 7.390000000e-07 V_low
+ 7.390010000e-07 V_low
+ 7.391000000e-07 V_low
+ 7.391010000e-07 V_low
+ 7.392000000e-07 V_low
+ 7.392010000e-07 V_low
+ 7.393000000e-07 V_low
+ 7.393010000e-07 V_low
+ 7.394000000e-07 V_low
+ 7.394010000e-07 V_low
+ 7.395000000e-07 V_low
+ 7.395010000e-07 V_low
+ 7.396000000e-07 V_low
+ 7.396010000e-07 V_low
+ 7.397000000e-07 V_low
+ 7.397010000e-07 V_low
+ 7.398000000e-07 V_low
+ 7.398010000e-07 V_low
+ 7.399000000e-07 V_low
+ 7.399010000e-07 V_low
+ 7.400000000e-07 V_low
+ 7.400010000e-07 V_low
+ 7.401000000e-07 V_low
+ 7.401010000e-07 V_low
+ 7.402000000e-07 V_low
+ 7.402010000e-07 V_low
+ 7.403000000e-07 V_low
+ 7.403010000e-07 V_low
+ 7.404000000e-07 V_low
+ 7.404010000e-07 V_low
+ 7.405000000e-07 V_low
+ 7.405010000e-07 V_low
+ 7.406000000e-07 V_low
+ 7.406010000e-07 V_low
+ 7.407000000e-07 V_low
+ 7.407010000e-07 V_low
+ 7.408000000e-07 V_low
+ 7.408010000e-07 V_low
+ 7.409000000e-07 V_low
+ 7.409010000e-07 V_low
+ 7.410000000e-07 V_low
+ 7.410010000e-07 V_low
+ 7.411000000e-07 V_low
+ 7.411010000e-07 V_low
+ 7.412000000e-07 V_low
+ 7.412010000e-07 V_low
+ 7.413000000e-07 V_low
+ 7.413010000e-07 V_low
+ 7.414000000e-07 V_low
+ 7.414010000e-07 V_low
+ 7.415000000e-07 V_low
+ 7.415010000e-07 V_low
+ 7.416000000e-07 V_low
+ 7.416010000e-07 V_low
+ 7.417000000e-07 V_low
+ 7.417010000e-07 V_low
+ 7.418000000e-07 V_low
+ 7.418010000e-07 V_low
+ 7.419000000e-07 V_low
+ 7.419010000e-07 V_low
+ 7.420000000e-07 V_low
+ 7.420010000e-07 V_low
+ 7.421000000e-07 V_low
+ 7.421010000e-07 V_low
+ 7.422000000e-07 V_low
+ 7.422010000e-07 V_low
+ 7.423000000e-07 V_low
+ 7.423010000e-07 V_low
+ 7.424000000e-07 V_low
+ 7.424010000e-07 V_low
+ 7.425000000e-07 V_low
+ 7.425010000e-07 V_low
+ 7.426000000e-07 V_low
+ 7.426010000e-07 V_low
+ 7.427000000e-07 V_low
+ 7.427010000e-07 V_low
+ 7.428000000e-07 V_low
+ 7.428010000e-07 V_low
+ 7.429000000e-07 V_low
+ 7.429010000e-07 V_hig
+ 7.430000000e-07 V_hig
+ 7.430010000e-07 V_hig
+ 7.431000000e-07 V_hig
+ 7.431010000e-07 V_hig
+ 7.432000000e-07 V_hig
+ 7.432010000e-07 V_hig
+ 7.433000000e-07 V_hig
+ 7.433010000e-07 V_hig
+ 7.434000000e-07 V_hig
+ 7.434010000e-07 V_hig
+ 7.435000000e-07 V_hig
+ 7.435010000e-07 V_hig
+ 7.436000000e-07 V_hig
+ 7.436010000e-07 V_hig
+ 7.437000000e-07 V_hig
+ 7.437010000e-07 V_hig
+ 7.438000000e-07 V_hig
+ 7.438010000e-07 V_hig
+ 7.439000000e-07 V_hig
+ 7.439010000e-07 V_low
+ 7.440000000e-07 V_low
+ 7.440010000e-07 V_low
+ 7.441000000e-07 V_low
+ 7.441010000e-07 V_low
+ 7.442000000e-07 V_low
+ 7.442010000e-07 V_low
+ 7.443000000e-07 V_low
+ 7.443010000e-07 V_low
+ 7.444000000e-07 V_low
+ 7.444010000e-07 V_low
+ 7.445000000e-07 V_low
+ 7.445010000e-07 V_low
+ 7.446000000e-07 V_low
+ 7.446010000e-07 V_low
+ 7.447000000e-07 V_low
+ 7.447010000e-07 V_low
+ 7.448000000e-07 V_low
+ 7.448010000e-07 V_low
+ 7.449000000e-07 V_low
+ 7.449010000e-07 V_low
+ 7.450000000e-07 V_low
+ 7.450010000e-07 V_low
+ 7.451000000e-07 V_low
+ 7.451010000e-07 V_low
+ 7.452000000e-07 V_low
+ 7.452010000e-07 V_low
+ 7.453000000e-07 V_low
+ 7.453010000e-07 V_low
+ 7.454000000e-07 V_low
+ 7.454010000e-07 V_low
+ 7.455000000e-07 V_low
+ 7.455010000e-07 V_low
+ 7.456000000e-07 V_low
+ 7.456010000e-07 V_low
+ 7.457000000e-07 V_low
+ 7.457010000e-07 V_low
+ 7.458000000e-07 V_low
+ 7.458010000e-07 V_low
+ 7.459000000e-07 V_low
+ 7.459010000e-07 V_low
+ 7.460000000e-07 V_low
+ 7.460010000e-07 V_low
+ 7.461000000e-07 V_low
+ 7.461010000e-07 V_low
+ 7.462000000e-07 V_low
+ 7.462010000e-07 V_low
+ 7.463000000e-07 V_low
+ 7.463010000e-07 V_low
+ 7.464000000e-07 V_low
+ 7.464010000e-07 V_low
+ 7.465000000e-07 V_low
+ 7.465010000e-07 V_low
+ 7.466000000e-07 V_low
+ 7.466010000e-07 V_low
+ 7.467000000e-07 V_low
+ 7.467010000e-07 V_low
+ 7.468000000e-07 V_low
+ 7.468010000e-07 V_low
+ 7.469000000e-07 V_low
+ 7.469010000e-07 V_low
+ 7.470000000e-07 V_low
+ 7.470010000e-07 V_low
+ 7.471000000e-07 V_low
+ 7.471010000e-07 V_low
+ 7.472000000e-07 V_low
+ 7.472010000e-07 V_low
+ 7.473000000e-07 V_low
+ 7.473010000e-07 V_low
+ 7.474000000e-07 V_low
+ 7.474010000e-07 V_low
+ 7.475000000e-07 V_low
+ 7.475010000e-07 V_low
+ 7.476000000e-07 V_low
+ 7.476010000e-07 V_low
+ 7.477000000e-07 V_low
+ 7.477010000e-07 V_low
+ 7.478000000e-07 V_low
+ 7.478010000e-07 V_low
+ 7.479000000e-07 V_low
+ 7.479010000e-07 V_hig
+ 7.480000000e-07 V_hig
+ 7.480010000e-07 V_hig
+ 7.481000000e-07 V_hig
+ 7.481010000e-07 V_hig
+ 7.482000000e-07 V_hig
+ 7.482010000e-07 V_hig
+ 7.483000000e-07 V_hig
+ 7.483010000e-07 V_hig
+ 7.484000000e-07 V_hig
+ 7.484010000e-07 V_hig
+ 7.485000000e-07 V_hig
+ 7.485010000e-07 V_hig
+ 7.486000000e-07 V_hig
+ 7.486010000e-07 V_hig
+ 7.487000000e-07 V_hig
+ 7.487010000e-07 V_hig
+ 7.488000000e-07 V_hig
+ 7.488010000e-07 V_hig
+ 7.489000000e-07 V_hig
+ 7.489010000e-07 V_hig
+ 7.490000000e-07 V_hig
+ 7.490010000e-07 V_hig
+ 7.491000000e-07 V_hig
+ 7.491010000e-07 V_hig
+ 7.492000000e-07 V_hig
+ 7.492010000e-07 V_hig
+ 7.493000000e-07 V_hig
+ 7.493010000e-07 V_hig
+ 7.494000000e-07 V_hig
+ 7.494010000e-07 V_hig
+ 7.495000000e-07 V_hig
+ 7.495010000e-07 V_hig
+ 7.496000000e-07 V_hig
+ 7.496010000e-07 V_hig
+ 7.497000000e-07 V_hig
+ 7.497010000e-07 V_hig
+ 7.498000000e-07 V_hig
+ 7.498010000e-07 V_hig
+ 7.499000000e-07 V_hig
+ 7.499010000e-07 V_low
+ 7.500000000e-07 V_low
+ 7.500010000e-07 V_low
+ 7.501000000e-07 V_low
+ 7.501010000e-07 V_low
+ 7.502000000e-07 V_low
+ 7.502010000e-07 V_low
+ 7.503000000e-07 V_low
+ 7.503010000e-07 V_low
+ 7.504000000e-07 V_low
+ 7.504010000e-07 V_low
+ 7.505000000e-07 V_low
+ 7.505010000e-07 V_low
+ 7.506000000e-07 V_low
+ 7.506010000e-07 V_low
+ 7.507000000e-07 V_low
+ 7.507010000e-07 V_low
+ 7.508000000e-07 V_low
+ 7.508010000e-07 V_low
+ 7.509000000e-07 V_low
+ 7.509010000e-07 V_hig
+ 7.510000000e-07 V_hig
+ 7.510010000e-07 V_hig
+ 7.511000000e-07 V_hig
+ 7.511010000e-07 V_hig
+ 7.512000000e-07 V_hig
+ 7.512010000e-07 V_hig
+ 7.513000000e-07 V_hig
+ 7.513010000e-07 V_hig
+ 7.514000000e-07 V_hig
+ 7.514010000e-07 V_hig
+ 7.515000000e-07 V_hig
+ 7.515010000e-07 V_hig
+ 7.516000000e-07 V_hig
+ 7.516010000e-07 V_hig
+ 7.517000000e-07 V_hig
+ 7.517010000e-07 V_hig
+ 7.518000000e-07 V_hig
+ 7.518010000e-07 V_hig
+ 7.519000000e-07 V_hig
+ 7.519010000e-07 V_hig
+ 7.520000000e-07 V_hig
+ 7.520010000e-07 V_hig
+ 7.521000000e-07 V_hig
+ 7.521010000e-07 V_hig
+ 7.522000000e-07 V_hig
+ 7.522010000e-07 V_hig
+ 7.523000000e-07 V_hig
+ 7.523010000e-07 V_hig
+ 7.524000000e-07 V_hig
+ 7.524010000e-07 V_hig
+ 7.525000000e-07 V_hig
+ 7.525010000e-07 V_hig
+ 7.526000000e-07 V_hig
+ 7.526010000e-07 V_hig
+ 7.527000000e-07 V_hig
+ 7.527010000e-07 V_hig
+ 7.528000000e-07 V_hig
+ 7.528010000e-07 V_hig
+ 7.529000000e-07 V_hig
+ 7.529010000e-07 V_hig
+ 7.530000000e-07 V_hig
+ 7.530010000e-07 V_hig
+ 7.531000000e-07 V_hig
+ 7.531010000e-07 V_hig
+ 7.532000000e-07 V_hig
+ 7.532010000e-07 V_hig
+ 7.533000000e-07 V_hig
+ 7.533010000e-07 V_hig
+ 7.534000000e-07 V_hig
+ 7.534010000e-07 V_hig
+ 7.535000000e-07 V_hig
+ 7.535010000e-07 V_hig
+ 7.536000000e-07 V_hig
+ 7.536010000e-07 V_hig
+ 7.537000000e-07 V_hig
+ 7.537010000e-07 V_hig
+ 7.538000000e-07 V_hig
+ 7.538010000e-07 V_hig
+ 7.539000000e-07 V_hig
+ 7.539010000e-07 V_low
+ 7.540000000e-07 V_low
+ 7.540010000e-07 V_low
+ 7.541000000e-07 V_low
+ 7.541010000e-07 V_low
+ 7.542000000e-07 V_low
+ 7.542010000e-07 V_low
+ 7.543000000e-07 V_low
+ 7.543010000e-07 V_low
+ 7.544000000e-07 V_low
+ 7.544010000e-07 V_low
+ 7.545000000e-07 V_low
+ 7.545010000e-07 V_low
+ 7.546000000e-07 V_low
+ 7.546010000e-07 V_low
+ 7.547000000e-07 V_low
+ 7.547010000e-07 V_low
+ 7.548000000e-07 V_low
+ 7.548010000e-07 V_low
+ 7.549000000e-07 V_low
+ 7.549010000e-07 V_hig
+ 7.550000000e-07 V_hig
+ 7.550010000e-07 V_hig
+ 7.551000000e-07 V_hig
+ 7.551010000e-07 V_hig
+ 7.552000000e-07 V_hig
+ 7.552010000e-07 V_hig
+ 7.553000000e-07 V_hig
+ 7.553010000e-07 V_hig
+ 7.554000000e-07 V_hig
+ 7.554010000e-07 V_hig
+ 7.555000000e-07 V_hig
+ 7.555010000e-07 V_hig
+ 7.556000000e-07 V_hig
+ 7.556010000e-07 V_hig
+ 7.557000000e-07 V_hig
+ 7.557010000e-07 V_hig
+ 7.558000000e-07 V_hig
+ 7.558010000e-07 V_hig
+ 7.559000000e-07 V_hig
+ 7.559010000e-07 V_hig
+ 7.560000000e-07 V_hig
+ 7.560010000e-07 V_hig
+ 7.561000000e-07 V_hig
+ 7.561010000e-07 V_hig
+ 7.562000000e-07 V_hig
+ 7.562010000e-07 V_hig
+ 7.563000000e-07 V_hig
+ 7.563010000e-07 V_hig
+ 7.564000000e-07 V_hig
+ 7.564010000e-07 V_hig
+ 7.565000000e-07 V_hig
+ 7.565010000e-07 V_hig
+ 7.566000000e-07 V_hig
+ 7.566010000e-07 V_hig
+ 7.567000000e-07 V_hig
+ 7.567010000e-07 V_hig
+ 7.568000000e-07 V_hig
+ 7.568010000e-07 V_hig
+ 7.569000000e-07 V_hig
+ 7.569010000e-07 V_hig
+ 7.570000000e-07 V_hig
+ 7.570010000e-07 V_hig
+ 7.571000000e-07 V_hig
+ 7.571010000e-07 V_hig
+ 7.572000000e-07 V_hig
+ 7.572010000e-07 V_hig
+ 7.573000000e-07 V_hig
+ 7.573010000e-07 V_hig
+ 7.574000000e-07 V_hig
+ 7.574010000e-07 V_hig
+ 7.575000000e-07 V_hig
+ 7.575010000e-07 V_hig
+ 7.576000000e-07 V_hig
+ 7.576010000e-07 V_hig
+ 7.577000000e-07 V_hig
+ 7.577010000e-07 V_hig
+ 7.578000000e-07 V_hig
+ 7.578010000e-07 V_hig
+ 7.579000000e-07 V_hig
+ 7.579010000e-07 V_low
+ 7.580000000e-07 V_low
+ 7.580010000e-07 V_low
+ 7.581000000e-07 V_low
+ 7.581010000e-07 V_low
+ 7.582000000e-07 V_low
+ 7.582010000e-07 V_low
+ 7.583000000e-07 V_low
+ 7.583010000e-07 V_low
+ 7.584000000e-07 V_low
+ 7.584010000e-07 V_low
+ 7.585000000e-07 V_low
+ 7.585010000e-07 V_low
+ 7.586000000e-07 V_low
+ 7.586010000e-07 V_low
+ 7.587000000e-07 V_low
+ 7.587010000e-07 V_low
+ 7.588000000e-07 V_low
+ 7.588010000e-07 V_low
+ 7.589000000e-07 V_low
+ 7.589010000e-07 V_low
+ 7.590000000e-07 V_low
+ 7.590010000e-07 V_low
+ 7.591000000e-07 V_low
+ 7.591010000e-07 V_low
+ 7.592000000e-07 V_low
+ 7.592010000e-07 V_low
+ 7.593000000e-07 V_low
+ 7.593010000e-07 V_low
+ 7.594000000e-07 V_low
+ 7.594010000e-07 V_low
+ 7.595000000e-07 V_low
+ 7.595010000e-07 V_low
+ 7.596000000e-07 V_low
+ 7.596010000e-07 V_low
+ 7.597000000e-07 V_low
+ 7.597010000e-07 V_low
+ 7.598000000e-07 V_low
+ 7.598010000e-07 V_low
+ 7.599000000e-07 V_low
+ 7.599010000e-07 V_low
+ 7.600000000e-07 V_low
+ 7.600010000e-07 V_low
+ 7.601000000e-07 V_low
+ 7.601010000e-07 V_low
+ 7.602000000e-07 V_low
+ 7.602010000e-07 V_low
+ 7.603000000e-07 V_low
+ 7.603010000e-07 V_low
+ 7.604000000e-07 V_low
+ 7.604010000e-07 V_low
+ 7.605000000e-07 V_low
+ 7.605010000e-07 V_low
+ 7.606000000e-07 V_low
+ 7.606010000e-07 V_low
+ 7.607000000e-07 V_low
+ 7.607010000e-07 V_low
+ 7.608000000e-07 V_low
+ 7.608010000e-07 V_low
+ 7.609000000e-07 V_low
+ 7.609010000e-07 V_hig
+ 7.610000000e-07 V_hig
+ 7.610010000e-07 V_hig
+ 7.611000000e-07 V_hig
+ 7.611010000e-07 V_hig
+ 7.612000000e-07 V_hig
+ 7.612010000e-07 V_hig
+ 7.613000000e-07 V_hig
+ 7.613010000e-07 V_hig
+ 7.614000000e-07 V_hig
+ 7.614010000e-07 V_hig
+ 7.615000000e-07 V_hig
+ 7.615010000e-07 V_hig
+ 7.616000000e-07 V_hig
+ 7.616010000e-07 V_hig
+ 7.617000000e-07 V_hig
+ 7.617010000e-07 V_hig
+ 7.618000000e-07 V_hig
+ 7.618010000e-07 V_hig
+ 7.619000000e-07 V_hig
+ 7.619010000e-07 V_hig
+ 7.620000000e-07 V_hig
+ 7.620010000e-07 V_hig
+ 7.621000000e-07 V_hig
+ 7.621010000e-07 V_hig
+ 7.622000000e-07 V_hig
+ 7.622010000e-07 V_hig
+ 7.623000000e-07 V_hig
+ 7.623010000e-07 V_hig
+ 7.624000000e-07 V_hig
+ 7.624010000e-07 V_hig
+ 7.625000000e-07 V_hig
+ 7.625010000e-07 V_hig
+ 7.626000000e-07 V_hig
+ 7.626010000e-07 V_hig
+ 7.627000000e-07 V_hig
+ 7.627010000e-07 V_hig
+ 7.628000000e-07 V_hig
+ 7.628010000e-07 V_hig
+ 7.629000000e-07 V_hig
+ 7.629010000e-07 V_low
+ 7.630000000e-07 V_low
+ 7.630010000e-07 V_low
+ 7.631000000e-07 V_low
+ 7.631010000e-07 V_low
+ 7.632000000e-07 V_low
+ 7.632010000e-07 V_low
+ 7.633000000e-07 V_low
+ 7.633010000e-07 V_low
+ 7.634000000e-07 V_low
+ 7.634010000e-07 V_low
+ 7.635000000e-07 V_low
+ 7.635010000e-07 V_low
+ 7.636000000e-07 V_low
+ 7.636010000e-07 V_low
+ 7.637000000e-07 V_low
+ 7.637010000e-07 V_low
+ 7.638000000e-07 V_low
+ 7.638010000e-07 V_low
+ 7.639000000e-07 V_low
+ 7.639010000e-07 V_low
+ 7.640000000e-07 V_low
+ 7.640010000e-07 V_low
+ 7.641000000e-07 V_low
+ 7.641010000e-07 V_low
+ 7.642000000e-07 V_low
+ 7.642010000e-07 V_low
+ 7.643000000e-07 V_low
+ 7.643010000e-07 V_low
+ 7.644000000e-07 V_low
+ 7.644010000e-07 V_low
+ 7.645000000e-07 V_low
+ 7.645010000e-07 V_low
+ 7.646000000e-07 V_low
+ 7.646010000e-07 V_low
+ 7.647000000e-07 V_low
+ 7.647010000e-07 V_low
+ 7.648000000e-07 V_low
+ 7.648010000e-07 V_low
+ 7.649000000e-07 V_low
+ 7.649010000e-07 V_hig
+ 7.650000000e-07 V_hig
+ 7.650010000e-07 V_hig
+ 7.651000000e-07 V_hig
+ 7.651010000e-07 V_hig
+ 7.652000000e-07 V_hig
+ 7.652010000e-07 V_hig
+ 7.653000000e-07 V_hig
+ 7.653010000e-07 V_hig
+ 7.654000000e-07 V_hig
+ 7.654010000e-07 V_hig
+ 7.655000000e-07 V_hig
+ 7.655010000e-07 V_hig
+ 7.656000000e-07 V_hig
+ 7.656010000e-07 V_hig
+ 7.657000000e-07 V_hig
+ 7.657010000e-07 V_hig
+ 7.658000000e-07 V_hig
+ 7.658010000e-07 V_hig
+ 7.659000000e-07 V_hig
+ 7.659010000e-07 V_low
+ 7.660000000e-07 V_low
+ 7.660010000e-07 V_low
+ 7.661000000e-07 V_low
+ 7.661010000e-07 V_low
+ 7.662000000e-07 V_low
+ 7.662010000e-07 V_low
+ 7.663000000e-07 V_low
+ 7.663010000e-07 V_low
+ 7.664000000e-07 V_low
+ 7.664010000e-07 V_low
+ 7.665000000e-07 V_low
+ 7.665010000e-07 V_low
+ 7.666000000e-07 V_low
+ 7.666010000e-07 V_low
+ 7.667000000e-07 V_low
+ 7.667010000e-07 V_low
+ 7.668000000e-07 V_low
+ 7.668010000e-07 V_low
+ 7.669000000e-07 V_low
+ 7.669010000e-07 V_low
+ 7.670000000e-07 V_low
+ 7.670010000e-07 V_low
+ 7.671000000e-07 V_low
+ 7.671010000e-07 V_low
+ 7.672000000e-07 V_low
+ 7.672010000e-07 V_low
+ 7.673000000e-07 V_low
+ 7.673010000e-07 V_low
+ 7.674000000e-07 V_low
+ 7.674010000e-07 V_low
+ 7.675000000e-07 V_low
+ 7.675010000e-07 V_low
+ 7.676000000e-07 V_low
+ 7.676010000e-07 V_low
+ 7.677000000e-07 V_low
+ 7.677010000e-07 V_low
+ 7.678000000e-07 V_low
+ 7.678010000e-07 V_low
+ 7.679000000e-07 V_low
+ 7.679010000e-07 V_hig
+ 7.680000000e-07 V_hig
+ 7.680010000e-07 V_hig
+ 7.681000000e-07 V_hig
+ 7.681010000e-07 V_hig
+ 7.682000000e-07 V_hig
+ 7.682010000e-07 V_hig
+ 7.683000000e-07 V_hig
+ 7.683010000e-07 V_hig
+ 7.684000000e-07 V_hig
+ 7.684010000e-07 V_hig
+ 7.685000000e-07 V_hig
+ 7.685010000e-07 V_hig
+ 7.686000000e-07 V_hig
+ 7.686010000e-07 V_hig
+ 7.687000000e-07 V_hig
+ 7.687010000e-07 V_hig
+ 7.688000000e-07 V_hig
+ 7.688010000e-07 V_hig
+ 7.689000000e-07 V_hig
+ 7.689010000e-07 V_hig
+ 7.690000000e-07 V_hig
+ 7.690010000e-07 V_hig
+ 7.691000000e-07 V_hig
+ 7.691010000e-07 V_hig
+ 7.692000000e-07 V_hig
+ 7.692010000e-07 V_hig
+ 7.693000000e-07 V_hig
+ 7.693010000e-07 V_hig
+ 7.694000000e-07 V_hig
+ 7.694010000e-07 V_hig
+ 7.695000000e-07 V_hig
+ 7.695010000e-07 V_hig
+ 7.696000000e-07 V_hig
+ 7.696010000e-07 V_hig
+ 7.697000000e-07 V_hig
+ 7.697010000e-07 V_hig
+ 7.698000000e-07 V_hig
+ 7.698010000e-07 V_hig
+ 7.699000000e-07 V_hig
+ 7.699010000e-07 V_hig
+ 7.700000000e-07 V_hig
+ 7.700010000e-07 V_hig
+ 7.701000000e-07 V_hig
+ 7.701010000e-07 V_hig
+ 7.702000000e-07 V_hig
+ 7.702010000e-07 V_hig
+ 7.703000000e-07 V_hig
+ 7.703010000e-07 V_hig
+ 7.704000000e-07 V_hig
+ 7.704010000e-07 V_hig
+ 7.705000000e-07 V_hig
+ 7.705010000e-07 V_hig
+ 7.706000000e-07 V_hig
+ 7.706010000e-07 V_hig
+ 7.707000000e-07 V_hig
+ 7.707010000e-07 V_hig
+ 7.708000000e-07 V_hig
+ 7.708010000e-07 V_hig
+ 7.709000000e-07 V_hig
+ 7.709010000e-07 V_hig
+ 7.710000000e-07 V_hig
+ 7.710010000e-07 V_hig
+ 7.711000000e-07 V_hig
+ 7.711010000e-07 V_hig
+ 7.712000000e-07 V_hig
+ 7.712010000e-07 V_hig
+ 7.713000000e-07 V_hig
+ 7.713010000e-07 V_hig
+ 7.714000000e-07 V_hig
+ 7.714010000e-07 V_hig
+ 7.715000000e-07 V_hig
+ 7.715010000e-07 V_hig
+ 7.716000000e-07 V_hig
+ 7.716010000e-07 V_hig
+ 7.717000000e-07 V_hig
+ 7.717010000e-07 V_hig
+ 7.718000000e-07 V_hig
+ 7.718010000e-07 V_hig
+ 7.719000000e-07 V_hig
+ 7.719010000e-07 V_hig
+ 7.720000000e-07 V_hig
+ 7.720010000e-07 V_hig
+ 7.721000000e-07 V_hig
+ 7.721010000e-07 V_hig
+ 7.722000000e-07 V_hig
+ 7.722010000e-07 V_hig
+ 7.723000000e-07 V_hig
+ 7.723010000e-07 V_hig
+ 7.724000000e-07 V_hig
+ 7.724010000e-07 V_hig
+ 7.725000000e-07 V_hig
+ 7.725010000e-07 V_hig
+ 7.726000000e-07 V_hig
+ 7.726010000e-07 V_hig
+ 7.727000000e-07 V_hig
+ 7.727010000e-07 V_hig
+ 7.728000000e-07 V_hig
+ 7.728010000e-07 V_hig
+ 7.729000000e-07 V_hig
+ 7.729010000e-07 V_hig
+ 7.730000000e-07 V_hig
+ 7.730010000e-07 V_hig
+ 7.731000000e-07 V_hig
+ 7.731010000e-07 V_hig
+ 7.732000000e-07 V_hig
+ 7.732010000e-07 V_hig
+ 7.733000000e-07 V_hig
+ 7.733010000e-07 V_hig
+ 7.734000000e-07 V_hig
+ 7.734010000e-07 V_hig
+ 7.735000000e-07 V_hig
+ 7.735010000e-07 V_hig
+ 7.736000000e-07 V_hig
+ 7.736010000e-07 V_hig
+ 7.737000000e-07 V_hig
+ 7.737010000e-07 V_hig
+ 7.738000000e-07 V_hig
+ 7.738010000e-07 V_hig
+ 7.739000000e-07 V_hig
+ 7.739010000e-07 V_low
+ 7.740000000e-07 V_low
+ 7.740010000e-07 V_low
+ 7.741000000e-07 V_low
+ 7.741010000e-07 V_low
+ 7.742000000e-07 V_low
+ 7.742010000e-07 V_low
+ 7.743000000e-07 V_low
+ 7.743010000e-07 V_low
+ 7.744000000e-07 V_low
+ 7.744010000e-07 V_low
+ 7.745000000e-07 V_low
+ 7.745010000e-07 V_low
+ 7.746000000e-07 V_low
+ 7.746010000e-07 V_low
+ 7.747000000e-07 V_low
+ 7.747010000e-07 V_low
+ 7.748000000e-07 V_low
+ 7.748010000e-07 V_low
+ 7.749000000e-07 V_low
+ 7.749010000e-07 V_hig
+ 7.750000000e-07 V_hig
+ 7.750010000e-07 V_hig
+ 7.751000000e-07 V_hig
+ 7.751010000e-07 V_hig
+ 7.752000000e-07 V_hig
+ 7.752010000e-07 V_hig
+ 7.753000000e-07 V_hig
+ 7.753010000e-07 V_hig
+ 7.754000000e-07 V_hig
+ 7.754010000e-07 V_hig
+ 7.755000000e-07 V_hig
+ 7.755010000e-07 V_hig
+ 7.756000000e-07 V_hig
+ 7.756010000e-07 V_hig
+ 7.757000000e-07 V_hig
+ 7.757010000e-07 V_hig
+ 7.758000000e-07 V_hig
+ 7.758010000e-07 V_hig
+ 7.759000000e-07 V_hig
+ 7.759010000e-07 V_hig
+ 7.760000000e-07 V_hig
+ 7.760010000e-07 V_hig
+ 7.761000000e-07 V_hig
+ 7.761010000e-07 V_hig
+ 7.762000000e-07 V_hig
+ 7.762010000e-07 V_hig
+ 7.763000000e-07 V_hig
+ 7.763010000e-07 V_hig
+ 7.764000000e-07 V_hig
+ 7.764010000e-07 V_hig
+ 7.765000000e-07 V_hig
+ 7.765010000e-07 V_hig
+ 7.766000000e-07 V_hig
+ 7.766010000e-07 V_hig
+ 7.767000000e-07 V_hig
+ 7.767010000e-07 V_hig
+ 7.768000000e-07 V_hig
+ 7.768010000e-07 V_hig
+ 7.769000000e-07 V_hig
+ 7.769010000e-07 V_low
+ 7.770000000e-07 V_low
+ 7.770010000e-07 V_low
+ 7.771000000e-07 V_low
+ 7.771010000e-07 V_low
+ 7.772000000e-07 V_low
+ 7.772010000e-07 V_low
+ 7.773000000e-07 V_low
+ 7.773010000e-07 V_low
+ 7.774000000e-07 V_low
+ 7.774010000e-07 V_low
+ 7.775000000e-07 V_low
+ 7.775010000e-07 V_low
+ 7.776000000e-07 V_low
+ 7.776010000e-07 V_low
+ 7.777000000e-07 V_low
+ 7.777010000e-07 V_low
+ 7.778000000e-07 V_low
+ 7.778010000e-07 V_low
+ 7.779000000e-07 V_low
+ 7.779010000e-07 V_low
+ 7.780000000e-07 V_low
+ 7.780010000e-07 V_low
+ 7.781000000e-07 V_low
+ 7.781010000e-07 V_low
+ 7.782000000e-07 V_low
+ 7.782010000e-07 V_low
+ 7.783000000e-07 V_low
+ 7.783010000e-07 V_low
+ 7.784000000e-07 V_low
+ 7.784010000e-07 V_low
+ 7.785000000e-07 V_low
+ 7.785010000e-07 V_low
+ 7.786000000e-07 V_low
+ 7.786010000e-07 V_low
+ 7.787000000e-07 V_low
+ 7.787010000e-07 V_low
+ 7.788000000e-07 V_low
+ 7.788010000e-07 V_low
+ 7.789000000e-07 V_low
+ 7.789010000e-07 V_low
+ 7.790000000e-07 V_low
+ 7.790010000e-07 V_low
+ 7.791000000e-07 V_low
+ 7.791010000e-07 V_low
+ 7.792000000e-07 V_low
+ 7.792010000e-07 V_low
+ 7.793000000e-07 V_low
+ 7.793010000e-07 V_low
+ 7.794000000e-07 V_low
+ 7.794010000e-07 V_low
+ 7.795000000e-07 V_low
+ 7.795010000e-07 V_low
+ 7.796000000e-07 V_low
+ 7.796010000e-07 V_low
+ 7.797000000e-07 V_low
+ 7.797010000e-07 V_low
+ 7.798000000e-07 V_low
+ 7.798010000e-07 V_low
+ 7.799000000e-07 V_low
+ 7.799010000e-07 V_low
+ 7.800000000e-07 V_low
+ 7.800010000e-07 V_low
+ 7.801000000e-07 V_low
+ 7.801010000e-07 V_low
+ 7.802000000e-07 V_low
+ 7.802010000e-07 V_low
+ 7.803000000e-07 V_low
+ 7.803010000e-07 V_low
+ 7.804000000e-07 V_low
+ 7.804010000e-07 V_low
+ 7.805000000e-07 V_low
+ 7.805010000e-07 V_low
+ 7.806000000e-07 V_low
+ 7.806010000e-07 V_low
+ 7.807000000e-07 V_low
+ 7.807010000e-07 V_low
+ 7.808000000e-07 V_low
+ 7.808010000e-07 V_low
+ 7.809000000e-07 V_low
+ 7.809010000e-07 V_low
+ 7.810000000e-07 V_low
+ 7.810010000e-07 V_low
+ 7.811000000e-07 V_low
+ 7.811010000e-07 V_low
+ 7.812000000e-07 V_low
+ 7.812010000e-07 V_low
+ 7.813000000e-07 V_low
+ 7.813010000e-07 V_low
+ 7.814000000e-07 V_low
+ 7.814010000e-07 V_low
+ 7.815000000e-07 V_low
+ 7.815010000e-07 V_low
+ 7.816000000e-07 V_low
+ 7.816010000e-07 V_low
+ 7.817000000e-07 V_low
+ 7.817010000e-07 V_low
+ 7.818000000e-07 V_low
+ 7.818010000e-07 V_low
+ 7.819000000e-07 V_low
+ 7.819010000e-07 V_hig
+ 7.820000000e-07 V_hig
+ 7.820010000e-07 V_hig
+ 7.821000000e-07 V_hig
+ 7.821010000e-07 V_hig
+ 7.822000000e-07 V_hig
+ 7.822010000e-07 V_hig
+ 7.823000000e-07 V_hig
+ 7.823010000e-07 V_hig
+ 7.824000000e-07 V_hig
+ 7.824010000e-07 V_hig
+ 7.825000000e-07 V_hig
+ 7.825010000e-07 V_hig
+ 7.826000000e-07 V_hig
+ 7.826010000e-07 V_hig
+ 7.827000000e-07 V_hig
+ 7.827010000e-07 V_hig
+ 7.828000000e-07 V_hig
+ 7.828010000e-07 V_hig
+ 7.829000000e-07 V_hig
+ 7.829010000e-07 V_hig
+ 7.830000000e-07 V_hig
+ 7.830010000e-07 V_hig
+ 7.831000000e-07 V_hig
+ 7.831010000e-07 V_hig
+ 7.832000000e-07 V_hig
+ 7.832010000e-07 V_hig
+ 7.833000000e-07 V_hig
+ 7.833010000e-07 V_hig
+ 7.834000000e-07 V_hig
+ 7.834010000e-07 V_hig
+ 7.835000000e-07 V_hig
+ 7.835010000e-07 V_hig
+ 7.836000000e-07 V_hig
+ 7.836010000e-07 V_hig
+ 7.837000000e-07 V_hig
+ 7.837010000e-07 V_hig
+ 7.838000000e-07 V_hig
+ 7.838010000e-07 V_hig
+ 7.839000000e-07 V_hig
+ 7.839010000e-07 V_hig
+ 7.840000000e-07 V_hig
+ 7.840010000e-07 V_hig
+ 7.841000000e-07 V_hig
+ 7.841010000e-07 V_hig
+ 7.842000000e-07 V_hig
+ 7.842010000e-07 V_hig
+ 7.843000000e-07 V_hig
+ 7.843010000e-07 V_hig
+ 7.844000000e-07 V_hig
+ 7.844010000e-07 V_hig
+ 7.845000000e-07 V_hig
+ 7.845010000e-07 V_hig
+ 7.846000000e-07 V_hig
+ 7.846010000e-07 V_hig
+ 7.847000000e-07 V_hig
+ 7.847010000e-07 V_hig
+ 7.848000000e-07 V_hig
+ 7.848010000e-07 V_hig
+ 7.849000000e-07 V_hig
+ 7.849010000e-07 V_hig
+ 7.850000000e-07 V_hig
+ 7.850010000e-07 V_hig
+ 7.851000000e-07 V_hig
+ 7.851010000e-07 V_hig
+ 7.852000000e-07 V_hig
+ 7.852010000e-07 V_hig
+ 7.853000000e-07 V_hig
+ 7.853010000e-07 V_hig
+ 7.854000000e-07 V_hig
+ 7.854010000e-07 V_hig
+ 7.855000000e-07 V_hig
+ 7.855010000e-07 V_hig
+ 7.856000000e-07 V_hig
+ 7.856010000e-07 V_hig
+ 7.857000000e-07 V_hig
+ 7.857010000e-07 V_hig
+ 7.858000000e-07 V_hig
+ 7.858010000e-07 V_hig
+ 7.859000000e-07 V_hig
+ 7.859010000e-07 V_low
+ 7.860000000e-07 V_low
+ 7.860010000e-07 V_low
+ 7.861000000e-07 V_low
+ 7.861010000e-07 V_low
+ 7.862000000e-07 V_low
+ 7.862010000e-07 V_low
+ 7.863000000e-07 V_low
+ 7.863010000e-07 V_low
+ 7.864000000e-07 V_low
+ 7.864010000e-07 V_low
+ 7.865000000e-07 V_low
+ 7.865010000e-07 V_low
+ 7.866000000e-07 V_low
+ 7.866010000e-07 V_low
+ 7.867000000e-07 V_low
+ 7.867010000e-07 V_low
+ 7.868000000e-07 V_low
+ 7.868010000e-07 V_low
+ 7.869000000e-07 V_low
+ 7.869010000e-07 V_hig
+ 7.870000000e-07 V_hig
+ 7.870010000e-07 V_hig
+ 7.871000000e-07 V_hig
+ 7.871010000e-07 V_hig
+ 7.872000000e-07 V_hig
+ 7.872010000e-07 V_hig
+ 7.873000000e-07 V_hig
+ 7.873010000e-07 V_hig
+ 7.874000000e-07 V_hig
+ 7.874010000e-07 V_hig
+ 7.875000000e-07 V_hig
+ 7.875010000e-07 V_hig
+ 7.876000000e-07 V_hig
+ 7.876010000e-07 V_hig
+ 7.877000000e-07 V_hig
+ 7.877010000e-07 V_hig
+ 7.878000000e-07 V_hig
+ 7.878010000e-07 V_hig
+ 7.879000000e-07 V_hig
+ 7.879010000e-07 V_low
+ 7.880000000e-07 V_low
+ 7.880010000e-07 V_low
+ 7.881000000e-07 V_low
+ 7.881010000e-07 V_low
+ 7.882000000e-07 V_low
+ 7.882010000e-07 V_low
+ 7.883000000e-07 V_low
+ 7.883010000e-07 V_low
+ 7.884000000e-07 V_low
+ 7.884010000e-07 V_low
+ 7.885000000e-07 V_low
+ 7.885010000e-07 V_low
+ 7.886000000e-07 V_low
+ 7.886010000e-07 V_low
+ 7.887000000e-07 V_low
+ 7.887010000e-07 V_low
+ 7.888000000e-07 V_low
+ 7.888010000e-07 V_low
+ 7.889000000e-07 V_low
+ 7.889010000e-07 V_hig
+ 7.890000000e-07 V_hig
+ 7.890010000e-07 V_hig
+ 7.891000000e-07 V_hig
+ 7.891010000e-07 V_hig
+ 7.892000000e-07 V_hig
+ 7.892010000e-07 V_hig
+ 7.893000000e-07 V_hig
+ 7.893010000e-07 V_hig
+ 7.894000000e-07 V_hig
+ 7.894010000e-07 V_hig
+ 7.895000000e-07 V_hig
+ 7.895010000e-07 V_hig
+ 7.896000000e-07 V_hig
+ 7.896010000e-07 V_hig
+ 7.897000000e-07 V_hig
+ 7.897010000e-07 V_hig
+ 7.898000000e-07 V_hig
+ 7.898010000e-07 V_hig
+ 7.899000000e-07 V_hig
+ 7.899010000e-07 V_hig
+ 7.900000000e-07 V_hig
+ 7.900010000e-07 V_hig
+ 7.901000000e-07 V_hig
+ 7.901010000e-07 V_hig
+ 7.902000000e-07 V_hig
+ 7.902010000e-07 V_hig
+ 7.903000000e-07 V_hig
+ 7.903010000e-07 V_hig
+ 7.904000000e-07 V_hig
+ 7.904010000e-07 V_hig
+ 7.905000000e-07 V_hig
+ 7.905010000e-07 V_hig
+ 7.906000000e-07 V_hig
+ 7.906010000e-07 V_hig
+ 7.907000000e-07 V_hig
+ 7.907010000e-07 V_hig
+ 7.908000000e-07 V_hig
+ 7.908010000e-07 V_hig
+ 7.909000000e-07 V_hig
+ 7.909010000e-07 V_hig
+ 7.910000000e-07 V_hig
+ 7.910010000e-07 V_hig
+ 7.911000000e-07 V_hig
+ 7.911010000e-07 V_hig
+ 7.912000000e-07 V_hig
+ 7.912010000e-07 V_hig
+ 7.913000000e-07 V_hig
+ 7.913010000e-07 V_hig
+ 7.914000000e-07 V_hig
+ 7.914010000e-07 V_hig
+ 7.915000000e-07 V_hig
+ 7.915010000e-07 V_hig
+ 7.916000000e-07 V_hig
+ 7.916010000e-07 V_hig
+ 7.917000000e-07 V_hig
+ 7.917010000e-07 V_hig
+ 7.918000000e-07 V_hig
+ 7.918010000e-07 V_hig
+ 7.919000000e-07 V_hig
+ 7.919010000e-07 V_low
+ 7.920000000e-07 V_low
+ 7.920010000e-07 V_low
+ 7.921000000e-07 V_low
+ 7.921010000e-07 V_low
+ 7.922000000e-07 V_low
+ 7.922010000e-07 V_low
+ 7.923000000e-07 V_low
+ 7.923010000e-07 V_low
+ 7.924000000e-07 V_low
+ 7.924010000e-07 V_low
+ 7.925000000e-07 V_low
+ 7.925010000e-07 V_low
+ 7.926000000e-07 V_low
+ 7.926010000e-07 V_low
+ 7.927000000e-07 V_low
+ 7.927010000e-07 V_low
+ 7.928000000e-07 V_low
+ 7.928010000e-07 V_low
+ 7.929000000e-07 V_low
+ 7.929010000e-07 V_hig
+ 7.930000000e-07 V_hig
+ 7.930010000e-07 V_hig
+ 7.931000000e-07 V_hig
+ 7.931010000e-07 V_hig
+ 7.932000000e-07 V_hig
+ 7.932010000e-07 V_hig
+ 7.933000000e-07 V_hig
+ 7.933010000e-07 V_hig
+ 7.934000000e-07 V_hig
+ 7.934010000e-07 V_hig
+ 7.935000000e-07 V_hig
+ 7.935010000e-07 V_hig
+ 7.936000000e-07 V_hig
+ 7.936010000e-07 V_hig
+ 7.937000000e-07 V_hig
+ 7.937010000e-07 V_hig
+ 7.938000000e-07 V_hig
+ 7.938010000e-07 V_hig
+ 7.939000000e-07 V_hig
+ 7.939010000e-07 V_low
+ 7.940000000e-07 V_low
+ 7.940010000e-07 V_low
+ 7.941000000e-07 V_low
+ 7.941010000e-07 V_low
+ 7.942000000e-07 V_low
+ 7.942010000e-07 V_low
+ 7.943000000e-07 V_low
+ 7.943010000e-07 V_low
+ 7.944000000e-07 V_low
+ 7.944010000e-07 V_low
+ 7.945000000e-07 V_low
+ 7.945010000e-07 V_low
+ 7.946000000e-07 V_low
+ 7.946010000e-07 V_low
+ 7.947000000e-07 V_low
+ 7.947010000e-07 V_low
+ 7.948000000e-07 V_low
+ 7.948010000e-07 V_low
+ 7.949000000e-07 V_low
+ 7.949010000e-07 V_hig
+ 7.950000000e-07 V_hig
+ 7.950010000e-07 V_hig
+ 7.951000000e-07 V_hig
+ 7.951010000e-07 V_hig
+ 7.952000000e-07 V_hig
+ 7.952010000e-07 V_hig
+ 7.953000000e-07 V_hig
+ 7.953010000e-07 V_hig
+ 7.954000000e-07 V_hig
+ 7.954010000e-07 V_hig
+ 7.955000000e-07 V_hig
+ 7.955010000e-07 V_hig
+ 7.956000000e-07 V_hig
+ 7.956010000e-07 V_hig
+ 7.957000000e-07 V_hig
+ 7.957010000e-07 V_hig
+ 7.958000000e-07 V_hig
+ 7.958010000e-07 V_hig
+ 7.959000000e-07 V_hig
+ 7.959010000e-07 V_hig
+ 7.960000000e-07 V_hig
+ 7.960010000e-07 V_hig
+ 7.961000000e-07 V_hig
+ 7.961010000e-07 V_hig
+ 7.962000000e-07 V_hig
+ 7.962010000e-07 V_hig
+ 7.963000000e-07 V_hig
+ 7.963010000e-07 V_hig
+ 7.964000000e-07 V_hig
+ 7.964010000e-07 V_hig
+ 7.965000000e-07 V_hig
+ 7.965010000e-07 V_hig
+ 7.966000000e-07 V_hig
+ 7.966010000e-07 V_hig
+ 7.967000000e-07 V_hig
+ 7.967010000e-07 V_hig
+ 7.968000000e-07 V_hig
+ 7.968010000e-07 V_hig
+ 7.969000000e-07 V_hig
+ 7.969010000e-07 V_hig
+ 7.970000000e-07 V_hig
+ 7.970010000e-07 V_hig
+ 7.971000000e-07 V_hig
+ 7.971010000e-07 V_hig
+ 7.972000000e-07 V_hig
+ 7.972010000e-07 V_hig
+ 7.973000000e-07 V_hig
+ 7.973010000e-07 V_hig
+ 7.974000000e-07 V_hig
+ 7.974010000e-07 V_hig
+ 7.975000000e-07 V_hig
+ 7.975010000e-07 V_hig
+ 7.976000000e-07 V_hig
+ 7.976010000e-07 V_hig
+ 7.977000000e-07 V_hig
+ 7.977010000e-07 V_hig
+ 7.978000000e-07 V_hig
+ 7.978010000e-07 V_hig
+ 7.979000000e-07 V_hig
+ 7.979010000e-07 V_low
+ 7.980000000e-07 V_low
+ 7.980010000e-07 V_low
+ 7.981000000e-07 V_low
+ 7.981010000e-07 V_low
+ 7.982000000e-07 V_low
+ 7.982010000e-07 V_low
+ 7.983000000e-07 V_low
+ 7.983010000e-07 V_low
+ 7.984000000e-07 V_low
+ 7.984010000e-07 V_low
+ 7.985000000e-07 V_low
+ 7.985010000e-07 V_low
+ 7.986000000e-07 V_low
+ 7.986010000e-07 V_low
+ 7.987000000e-07 V_low
+ 7.987010000e-07 V_low
+ 7.988000000e-07 V_low
+ 7.988010000e-07 V_low
+ 7.989000000e-07 V_low
+ 7.989010000e-07 V_low
+ 7.990000000e-07 V_low
+ 7.990010000e-07 V_low
+ 7.991000000e-07 V_low
+ 7.991010000e-07 V_low
+ 7.992000000e-07 V_low
+ 7.992010000e-07 V_low
+ 7.993000000e-07 V_low
+ 7.993010000e-07 V_low
+ 7.994000000e-07 V_low
+ 7.994010000e-07 V_low
+ 7.995000000e-07 V_low
+ 7.995010000e-07 V_low
+ 7.996000000e-07 V_low
+ 7.996010000e-07 V_low
+ 7.997000000e-07 V_low
+ 7.997010000e-07 V_low
+ 7.998000000e-07 V_low
+ 7.998010000e-07 V_low
+ 7.999000000e-07 V_low
+ 7.999010000e-07 V_low
+ 8.000000000e-07 V_low
+ 8.000010000e-07 V_low
+ 8.001000000e-07 V_low
+ 8.001010000e-07 V_low
+ 8.002000000e-07 V_low
+ 8.002010000e-07 V_low
+ 8.003000000e-07 V_low
+ 8.003010000e-07 V_low
+ 8.004000000e-07 V_low
+ 8.004010000e-07 V_low
+ 8.005000000e-07 V_low
+ 8.005010000e-07 V_low
+ 8.006000000e-07 V_low
+ 8.006010000e-07 V_low
+ 8.007000000e-07 V_low
+ 8.007010000e-07 V_low
+ 8.008000000e-07 V_low
+ 8.008010000e-07 V_low
+ 8.009000000e-07 V_low
+ 8.009010000e-07 V_hig
+ 8.010000000e-07 V_hig
+ 8.010010000e-07 V_hig
+ 8.011000000e-07 V_hig
+ 8.011010000e-07 V_hig
+ 8.012000000e-07 V_hig
+ 8.012010000e-07 V_hig
+ 8.013000000e-07 V_hig
+ 8.013010000e-07 V_hig
+ 8.014000000e-07 V_hig
+ 8.014010000e-07 V_hig
+ 8.015000000e-07 V_hig
+ 8.015010000e-07 V_hig
+ 8.016000000e-07 V_hig
+ 8.016010000e-07 V_hig
+ 8.017000000e-07 V_hig
+ 8.017010000e-07 V_hig
+ 8.018000000e-07 V_hig
+ 8.018010000e-07 V_hig
+ 8.019000000e-07 V_hig
+ 8.019010000e-07 V_hig
+ 8.020000000e-07 V_hig
+ 8.020010000e-07 V_hig
+ 8.021000000e-07 V_hig
+ 8.021010000e-07 V_hig
+ 8.022000000e-07 V_hig
+ 8.022010000e-07 V_hig
+ 8.023000000e-07 V_hig
+ 8.023010000e-07 V_hig
+ 8.024000000e-07 V_hig
+ 8.024010000e-07 V_hig
+ 8.025000000e-07 V_hig
+ 8.025010000e-07 V_hig
+ 8.026000000e-07 V_hig
+ 8.026010000e-07 V_hig
+ 8.027000000e-07 V_hig
+ 8.027010000e-07 V_hig
+ 8.028000000e-07 V_hig
+ 8.028010000e-07 V_hig
+ 8.029000000e-07 V_hig
+ 8.029010000e-07 V_low
+ 8.030000000e-07 V_low
+ 8.030010000e-07 V_low
+ 8.031000000e-07 V_low
+ 8.031010000e-07 V_low
+ 8.032000000e-07 V_low
+ 8.032010000e-07 V_low
+ 8.033000000e-07 V_low
+ 8.033010000e-07 V_low
+ 8.034000000e-07 V_low
+ 8.034010000e-07 V_low
+ 8.035000000e-07 V_low
+ 8.035010000e-07 V_low
+ 8.036000000e-07 V_low
+ 8.036010000e-07 V_low
+ 8.037000000e-07 V_low
+ 8.037010000e-07 V_low
+ 8.038000000e-07 V_low
+ 8.038010000e-07 V_low
+ 8.039000000e-07 V_low
+ 8.039010000e-07 V_low
+ 8.040000000e-07 V_low
+ 8.040010000e-07 V_low
+ 8.041000000e-07 V_low
+ 8.041010000e-07 V_low
+ 8.042000000e-07 V_low
+ 8.042010000e-07 V_low
+ 8.043000000e-07 V_low
+ 8.043010000e-07 V_low
+ 8.044000000e-07 V_low
+ 8.044010000e-07 V_low
+ 8.045000000e-07 V_low
+ 8.045010000e-07 V_low
+ 8.046000000e-07 V_low
+ 8.046010000e-07 V_low
+ 8.047000000e-07 V_low
+ 8.047010000e-07 V_low
+ 8.048000000e-07 V_low
+ 8.048010000e-07 V_low
+ 8.049000000e-07 V_low
+ 8.049010000e-07 V_low
+ 8.050000000e-07 V_low
+ 8.050010000e-07 V_low
+ 8.051000000e-07 V_low
+ 8.051010000e-07 V_low
+ 8.052000000e-07 V_low
+ 8.052010000e-07 V_low
+ 8.053000000e-07 V_low
+ 8.053010000e-07 V_low
+ 8.054000000e-07 V_low
+ 8.054010000e-07 V_low
+ 8.055000000e-07 V_low
+ 8.055010000e-07 V_low
+ 8.056000000e-07 V_low
+ 8.056010000e-07 V_low
+ 8.057000000e-07 V_low
+ 8.057010000e-07 V_low
+ 8.058000000e-07 V_low
+ 8.058010000e-07 V_low
+ 8.059000000e-07 V_low
+ 8.059010000e-07 V_low
+ 8.060000000e-07 V_low
+ 8.060010000e-07 V_low
+ 8.061000000e-07 V_low
+ 8.061010000e-07 V_low
+ 8.062000000e-07 V_low
+ 8.062010000e-07 V_low
+ 8.063000000e-07 V_low
+ 8.063010000e-07 V_low
+ 8.064000000e-07 V_low
+ 8.064010000e-07 V_low
+ 8.065000000e-07 V_low
+ 8.065010000e-07 V_low
+ 8.066000000e-07 V_low
+ 8.066010000e-07 V_low
+ 8.067000000e-07 V_low
+ 8.067010000e-07 V_low
+ 8.068000000e-07 V_low
+ 8.068010000e-07 V_low
+ 8.069000000e-07 V_low
+ 8.069010000e-07 V_hig
+ 8.070000000e-07 V_hig
+ 8.070010000e-07 V_hig
+ 8.071000000e-07 V_hig
+ 8.071010000e-07 V_hig
+ 8.072000000e-07 V_hig
+ 8.072010000e-07 V_hig
+ 8.073000000e-07 V_hig
+ 8.073010000e-07 V_hig
+ 8.074000000e-07 V_hig
+ 8.074010000e-07 V_hig
+ 8.075000000e-07 V_hig
+ 8.075010000e-07 V_hig
+ 8.076000000e-07 V_hig
+ 8.076010000e-07 V_hig
+ 8.077000000e-07 V_hig
+ 8.077010000e-07 V_hig
+ 8.078000000e-07 V_hig
+ 8.078010000e-07 V_hig
+ 8.079000000e-07 V_hig
+ 8.079010000e-07 V_hig
+ 8.080000000e-07 V_hig
+ 8.080010000e-07 V_hig
+ 8.081000000e-07 V_hig
+ 8.081010000e-07 V_hig
+ 8.082000000e-07 V_hig
+ 8.082010000e-07 V_hig
+ 8.083000000e-07 V_hig
+ 8.083010000e-07 V_hig
+ 8.084000000e-07 V_hig
+ 8.084010000e-07 V_hig
+ 8.085000000e-07 V_hig
+ 8.085010000e-07 V_hig
+ 8.086000000e-07 V_hig
+ 8.086010000e-07 V_hig
+ 8.087000000e-07 V_hig
+ 8.087010000e-07 V_hig
+ 8.088000000e-07 V_hig
+ 8.088010000e-07 V_hig
+ 8.089000000e-07 V_hig
+ 8.089010000e-07 V_low
+ 8.090000000e-07 V_low
+ 8.090010000e-07 V_low
+ 8.091000000e-07 V_low
+ 8.091010000e-07 V_low
+ 8.092000000e-07 V_low
+ 8.092010000e-07 V_low
+ 8.093000000e-07 V_low
+ 8.093010000e-07 V_low
+ 8.094000000e-07 V_low
+ 8.094010000e-07 V_low
+ 8.095000000e-07 V_low
+ 8.095010000e-07 V_low
+ 8.096000000e-07 V_low
+ 8.096010000e-07 V_low
+ 8.097000000e-07 V_low
+ 8.097010000e-07 V_low
+ 8.098000000e-07 V_low
+ 8.098010000e-07 V_low
+ 8.099000000e-07 V_low
+ 8.099010000e-07 V_low
+ 8.100000000e-07 V_low
+ 8.100010000e-07 V_low
+ 8.101000000e-07 V_low
+ 8.101010000e-07 V_low
+ 8.102000000e-07 V_low
+ 8.102010000e-07 V_low
+ 8.103000000e-07 V_low
+ 8.103010000e-07 V_low
+ 8.104000000e-07 V_low
+ 8.104010000e-07 V_low
+ 8.105000000e-07 V_low
+ 8.105010000e-07 V_low
+ 8.106000000e-07 V_low
+ 8.106010000e-07 V_low
+ 8.107000000e-07 V_low
+ 8.107010000e-07 V_low
+ 8.108000000e-07 V_low
+ 8.108010000e-07 V_low
+ 8.109000000e-07 V_low
+ 8.109010000e-07 V_low
+ 8.110000000e-07 V_low
+ 8.110010000e-07 V_low
+ 8.111000000e-07 V_low
+ 8.111010000e-07 V_low
+ 8.112000000e-07 V_low
+ 8.112010000e-07 V_low
+ 8.113000000e-07 V_low
+ 8.113010000e-07 V_low
+ 8.114000000e-07 V_low
+ 8.114010000e-07 V_low
+ 8.115000000e-07 V_low
+ 8.115010000e-07 V_low
+ 8.116000000e-07 V_low
+ 8.116010000e-07 V_low
+ 8.117000000e-07 V_low
+ 8.117010000e-07 V_low
+ 8.118000000e-07 V_low
+ 8.118010000e-07 V_low
+ 8.119000000e-07 V_low
+ 8.119010000e-07 V_hig
+ 8.120000000e-07 V_hig
+ 8.120010000e-07 V_hig
+ 8.121000000e-07 V_hig
+ 8.121010000e-07 V_hig
+ 8.122000000e-07 V_hig
+ 8.122010000e-07 V_hig
+ 8.123000000e-07 V_hig
+ 8.123010000e-07 V_hig
+ 8.124000000e-07 V_hig
+ 8.124010000e-07 V_hig
+ 8.125000000e-07 V_hig
+ 8.125010000e-07 V_hig
+ 8.126000000e-07 V_hig
+ 8.126010000e-07 V_hig
+ 8.127000000e-07 V_hig
+ 8.127010000e-07 V_hig
+ 8.128000000e-07 V_hig
+ 8.128010000e-07 V_hig
+ 8.129000000e-07 V_hig
+ 8.129010000e-07 V_low
+ 8.130000000e-07 V_low
+ 8.130010000e-07 V_low
+ 8.131000000e-07 V_low
+ 8.131010000e-07 V_low
+ 8.132000000e-07 V_low
+ 8.132010000e-07 V_low
+ 8.133000000e-07 V_low
+ 8.133010000e-07 V_low
+ 8.134000000e-07 V_low
+ 8.134010000e-07 V_low
+ 8.135000000e-07 V_low
+ 8.135010000e-07 V_low
+ 8.136000000e-07 V_low
+ 8.136010000e-07 V_low
+ 8.137000000e-07 V_low
+ 8.137010000e-07 V_low
+ 8.138000000e-07 V_low
+ 8.138010000e-07 V_low
+ 8.139000000e-07 V_low
+ 8.139010000e-07 V_low
+ 8.140000000e-07 V_low
+ 8.140010000e-07 V_low
+ 8.141000000e-07 V_low
+ 8.141010000e-07 V_low
+ 8.142000000e-07 V_low
+ 8.142010000e-07 V_low
+ 8.143000000e-07 V_low
+ 8.143010000e-07 V_low
+ 8.144000000e-07 V_low
+ 8.144010000e-07 V_low
+ 8.145000000e-07 V_low
+ 8.145010000e-07 V_low
+ 8.146000000e-07 V_low
+ 8.146010000e-07 V_low
+ 8.147000000e-07 V_low
+ 8.147010000e-07 V_low
+ 8.148000000e-07 V_low
+ 8.148010000e-07 V_low
+ 8.149000000e-07 V_low
+ 8.149010000e-07 V_low
+ 8.150000000e-07 V_low
+ 8.150010000e-07 V_low
+ 8.151000000e-07 V_low
+ 8.151010000e-07 V_low
+ 8.152000000e-07 V_low
+ 8.152010000e-07 V_low
+ 8.153000000e-07 V_low
+ 8.153010000e-07 V_low
+ 8.154000000e-07 V_low
+ 8.154010000e-07 V_low
+ 8.155000000e-07 V_low
+ 8.155010000e-07 V_low
+ 8.156000000e-07 V_low
+ 8.156010000e-07 V_low
+ 8.157000000e-07 V_low
+ 8.157010000e-07 V_low
+ 8.158000000e-07 V_low
+ 8.158010000e-07 V_low
+ 8.159000000e-07 V_low
+ 8.159010000e-07 V_low
+ 8.160000000e-07 V_low
+ 8.160010000e-07 V_low
+ 8.161000000e-07 V_low
+ 8.161010000e-07 V_low
+ 8.162000000e-07 V_low
+ 8.162010000e-07 V_low
+ 8.163000000e-07 V_low
+ 8.163010000e-07 V_low
+ 8.164000000e-07 V_low
+ 8.164010000e-07 V_low
+ 8.165000000e-07 V_low
+ 8.165010000e-07 V_low
+ 8.166000000e-07 V_low
+ 8.166010000e-07 V_low
+ 8.167000000e-07 V_low
+ 8.167010000e-07 V_low
+ 8.168000000e-07 V_low
+ 8.168010000e-07 V_low
+ 8.169000000e-07 V_low
+ 8.169010000e-07 V_low
+ 8.170000000e-07 V_low
+ 8.170010000e-07 V_low
+ 8.171000000e-07 V_low
+ 8.171010000e-07 V_low
+ 8.172000000e-07 V_low
+ 8.172010000e-07 V_low
+ 8.173000000e-07 V_low
+ 8.173010000e-07 V_low
+ 8.174000000e-07 V_low
+ 8.174010000e-07 V_low
+ 8.175000000e-07 V_low
+ 8.175010000e-07 V_low
+ 8.176000000e-07 V_low
+ 8.176010000e-07 V_low
+ 8.177000000e-07 V_low
+ 8.177010000e-07 V_low
+ 8.178000000e-07 V_low
+ 8.178010000e-07 V_low
+ 8.179000000e-07 V_low
+ 8.179010000e-07 V_low
+ 8.180000000e-07 V_low
+ 8.180010000e-07 V_low
+ 8.181000000e-07 V_low
+ 8.181010000e-07 V_low
+ 8.182000000e-07 V_low
+ 8.182010000e-07 V_low
+ 8.183000000e-07 V_low
+ 8.183010000e-07 V_low
+ 8.184000000e-07 V_low
+ 8.184010000e-07 V_low
+ 8.185000000e-07 V_low
+ 8.185010000e-07 V_low
+ 8.186000000e-07 V_low
+ 8.186010000e-07 V_low
+ 8.187000000e-07 V_low
+ 8.187010000e-07 V_low
+ 8.188000000e-07 V_low
+ 8.188010000e-07 V_low
+ 8.189000000e-07 V_low
+ 8.189010000e-07 V_hig
+ 8.190000000e-07 V_hig
+ 8.190010000e-07 V_hig
+ 8.191000000e-07 V_hig
+ 8.191010000e-07 V_hig
+ 8.192000000e-07 V_hig
+ 8.192010000e-07 V_hig
+ 8.193000000e-07 V_hig
+ 8.193010000e-07 V_hig
+ 8.194000000e-07 V_hig
+ 8.194010000e-07 V_hig
+ 8.195000000e-07 V_hig
+ 8.195010000e-07 V_hig
+ 8.196000000e-07 V_hig
+ 8.196010000e-07 V_hig
+ 8.197000000e-07 V_hig
+ 8.197010000e-07 V_hig
+ 8.198000000e-07 V_hig
+ 8.198010000e-07 V_hig
+ 8.199000000e-07 V_hig
+ 8.199010000e-07 V_low
+ 8.200000000e-07 V_low
+ 8.200010000e-07 V_low
+ 8.201000000e-07 V_low
+ 8.201010000e-07 V_low
+ 8.202000000e-07 V_low
+ 8.202010000e-07 V_low
+ 8.203000000e-07 V_low
+ 8.203010000e-07 V_low
+ 8.204000000e-07 V_low
+ 8.204010000e-07 V_low
+ 8.205000000e-07 V_low
+ 8.205010000e-07 V_low
+ 8.206000000e-07 V_low
+ 8.206010000e-07 V_low
+ 8.207000000e-07 V_low
+ 8.207010000e-07 V_low
+ 8.208000000e-07 V_low
+ 8.208010000e-07 V_low
+ 8.209000000e-07 V_low
+ 8.209010000e-07 V_hig
+ 8.210000000e-07 V_hig
+ 8.210010000e-07 V_hig
+ 8.211000000e-07 V_hig
+ 8.211010000e-07 V_hig
+ 8.212000000e-07 V_hig
+ 8.212010000e-07 V_hig
+ 8.213000000e-07 V_hig
+ 8.213010000e-07 V_hig
+ 8.214000000e-07 V_hig
+ 8.214010000e-07 V_hig
+ 8.215000000e-07 V_hig
+ 8.215010000e-07 V_hig
+ 8.216000000e-07 V_hig
+ 8.216010000e-07 V_hig
+ 8.217000000e-07 V_hig
+ 8.217010000e-07 V_hig
+ 8.218000000e-07 V_hig
+ 8.218010000e-07 V_hig
+ 8.219000000e-07 V_hig
+ 8.219010000e-07 V_low
+ 8.220000000e-07 V_low
+ 8.220010000e-07 V_low
+ 8.221000000e-07 V_low
+ 8.221010000e-07 V_low
+ 8.222000000e-07 V_low
+ 8.222010000e-07 V_low
+ 8.223000000e-07 V_low
+ 8.223010000e-07 V_low
+ 8.224000000e-07 V_low
+ 8.224010000e-07 V_low
+ 8.225000000e-07 V_low
+ 8.225010000e-07 V_low
+ 8.226000000e-07 V_low
+ 8.226010000e-07 V_low
+ 8.227000000e-07 V_low
+ 8.227010000e-07 V_low
+ 8.228000000e-07 V_low
+ 8.228010000e-07 V_low
+ 8.229000000e-07 V_low
+ 8.229010000e-07 V_low
+ 8.230000000e-07 V_low
+ 8.230010000e-07 V_low
+ 8.231000000e-07 V_low
+ 8.231010000e-07 V_low
+ 8.232000000e-07 V_low
+ 8.232010000e-07 V_low
+ 8.233000000e-07 V_low
+ 8.233010000e-07 V_low
+ 8.234000000e-07 V_low
+ 8.234010000e-07 V_low
+ 8.235000000e-07 V_low
+ 8.235010000e-07 V_low
+ 8.236000000e-07 V_low
+ 8.236010000e-07 V_low
+ 8.237000000e-07 V_low
+ 8.237010000e-07 V_low
+ 8.238000000e-07 V_low
+ 8.238010000e-07 V_low
+ 8.239000000e-07 V_low
+ 8.239010000e-07 V_hig
+ 8.240000000e-07 V_hig
+ 8.240010000e-07 V_hig
+ 8.241000000e-07 V_hig
+ 8.241010000e-07 V_hig
+ 8.242000000e-07 V_hig
+ 8.242010000e-07 V_hig
+ 8.243000000e-07 V_hig
+ 8.243010000e-07 V_hig
+ 8.244000000e-07 V_hig
+ 8.244010000e-07 V_hig
+ 8.245000000e-07 V_hig
+ 8.245010000e-07 V_hig
+ 8.246000000e-07 V_hig
+ 8.246010000e-07 V_hig
+ 8.247000000e-07 V_hig
+ 8.247010000e-07 V_hig
+ 8.248000000e-07 V_hig
+ 8.248010000e-07 V_hig
+ 8.249000000e-07 V_hig
+ 8.249010000e-07 V_hig
+ 8.250000000e-07 V_hig
+ 8.250010000e-07 V_hig
+ 8.251000000e-07 V_hig
+ 8.251010000e-07 V_hig
+ 8.252000000e-07 V_hig
+ 8.252010000e-07 V_hig
+ 8.253000000e-07 V_hig
+ 8.253010000e-07 V_hig
+ 8.254000000e-07 V_hig
+ 8.254010000e-07 V_hig
+ 8.255000000e-07 V_hig
+ 8.255010000e-07 V_hig
+ 8.256000000e-07 V_hig
+ 8.256010000e-07 V_hig
+ 8.257000000e-07 V_hig
+ 8.257010000e-07 V_hig
+ 8.258000000e-07 V_hig
+ 8.258010000e-07 V_hig
+ 8.259000000e-07 V_hig
+ 8.259010000e-07 V_low
+ 8.260000000e-07 V_low
+ 8.260010000e-07 V_low
+ 8.261000000e-07 V_low
+ 8.261010000e-07 V_low
+ 8.262000000e-07 V_low
+ 8.262010000e-07 V_low
+ 8.263000000e-07 V_low
+ 8.263010000e-07 V_low
+ 8.264000000e-07 V_low
+ 8.264010000e-07 V_low
+ 8.265000000e-07 V_low
+ 8.265010000e-07 V_low
+ 8.266000000e-07 V_low
+ 8.266010000e-07 V_low
+ 8.267000000e-07 V_low
+ 8.267010000e-07 V_low
+ 8.268000000e-07 V_low
+ 8.268010000e-07 V_low
+ 8.269000000e-07 V_low
+ 8.269010000e-07 V_hig
+ 8.270000000e-07 V_hig
+ 8.270010000e-07 V_hig
+ 8.271000000e-07 V_hig
+ 8.271010000e-07 V_hig
+ 8.272000000e-07 V_hig
+ 8.272010000e-07 V_hig
+ 8.273000000e-07 V_hig
+ 8.273010000e-07 V_hig
+ 8.274000000e-07 V_hig
+ 8.274010000e-07 V_hig
+ 8.275000000e-07 V_hig
+ 8.275010000e-07 V_hig
+ 8.276000000e-07 V_hig
+ 8.276010000e-07 V_hig
+ 8.277000000e-07 V_hig
+ 8.277010000e-07 V_hig
+ 8.278000000e-07 V_hig
+ 8.278010000e-07 V_hig
+ 8.279000000e-07 V_hig
+ 8.279010000e-07 V_low
+ 8.280000000e-07 V_low
+ 8.280010000e-07 V_low
+ 8.281000000e-07 V_low
+ 8.281010000e-07 V_low
+ 8.282000000e-07 V_low
+ 8.282010000e-07 V_low
+ 8.283000000e-07 V_low
+ 8.283010000e-07 V_low
+ 8.284000000e-07 V_low
+ 8.284010000e-07 V_low
+ 8.285000000e-07 V_low
+ 8.285010000e-07 V_low
+ 8.286000000e-07 V_low
+ 8.286010000e-07 V_low
+ 8.287000000e-07 V_low
+ 8.287010000e-07 V_low
+ 8.288000000e-07 V_low
+ 8.288010000e-07 V_low
+ 8.289000000e-07 V_low
+ 8.289010000e-07 V_low
+ 8.290000000e-07 V_low
+ 8.290010000e-07 V_low
+ 8.291000000e-07 V_low
+ 8.291010000e-07 V_low
+ 8.292000000e-07 V_low
+ 8.292010000e-07 V_low
+ 8.293000000e-07 V_low
+ 8.293010000e-07 V_low
+ 8.294000000e-07 V_low
+ 8.294010000e-07 V_low
+ 8.295000000e-07 V_low
+ 8.295010000e-07 V_low
+ 8.296000000e-07 V_low
+ 8.296010000e-07 V_low
+ 8.297000000e-07 V_low
+ 8.297010000e-07 V_low
+ 8.298000000e-07 V_low
+ 8.298010000e-07 V_low
+ 8.299000000e-07 V_low
+ 8.299010000e-07 V_hig
+ 8.300000000e-07 V_hig
+ 8.300010000e-07 V_hig
+ 8.301000000e-07 V_hig
+ 8.301010000e-07 V_hig
+ 8.302000000e-07 V_hig
+ 8.302010000e-07 V_hig
+ 8.303000000e-07 V_hig
+ 8.303010000e-07 V_hig
+ 8.304000000e-07 V_hig
+ 8.304010000e-07 V_hig
+ 8.305000000e-07 V_hig
+ 8.305010000e-07 V_hig
+ 8.306000000e-07 V_hig
+ 8.306010000e-07 V_hig
+ 8.307000000e-07 V_hig
+ 8.307010000e-07 V_hig
+ 8.308000000e-07 V_hig
+ 8.308010000e-07 V_hig
+ 8.309000000e-07 V_hig
+ 8.309010000e-07 V_low
+ 8.310000000e-07 V_low
+ 8.310010000e-07 V_low
+ 8.311000000e-07 V_low
+ 8.311010000e-07 V_low
+ 8.312000000e-07 V_low
+ 8.312010000e-07 V_low
+ 8.313000000e-07 V_low
+ 8.313010000e-07 V_low
+ 8.314000000e-07 V_low
+ 8.314010000e-07 V_low
+ 8.315000000e-07 V_low
+ 8.315010000e-07 V_low
+ 8.316000000e-07 V_low
+ 8.316010000e-07 V_low
+ 8.317000000e-07 V_low
+ 8.317010000e-07 V_low
+ 8.318000000e-07 V_low
+ 8.318010000e-07 V_low
+ 8.319000000e-07 V_low
+ 8.319010000e-07 V_low
+ 8.320000000e-07 V_low
+ 8.320010000e-07 V_low
+ 8.321000000e-07 V_low
+ 8.321010000e-07 V_low
+ 8.322000000e-07 V_low
+ 8.322010000e-07 V_low
+ 8.323000000e-07 V_low
+ 8.323010000e-07 V_low
+ 8.324000000e-07 V_low
+ 8.324010000e-07 V_low
+ 8.325000000e-07 V_low
+ 8.325010000e-07 V_low
+ 8.326000000e-07 V_low
+ 8.326010000e-07 V_low
+ 8.327000000e-07 V_low
+ 8.327010000e-07 V_low
+ 8.328000000e-07 V_low
+ 8.328010000e-07 V_low
+ 8.329000000e-07 V_low
+ 8.329010000e-07 V_low
+ 8.330000000e-07 V_low
+ 8.330010000e-07 V_low
+ 8.331000000e-07 V_low
+ 8.331010000e-07 V_low
+ 8.332000000e-07 V_low
+ 8.332010000e-07 V_low
+ 8.333000000e-07 V_low
+ 8.333010000e-07 V_low
+ 8.334000000e-07 V_low
+ 8.334010000e-07 V_low
+ 8.335000000e-07 V_low
+ 8.335010000e-07 V_low
+ 8.336000000e-07 V_low
+ 8.336010000e-07 V_low
+ 8.337000000e-07 V_low
+ 8.337010000e-07 V_low
+ 8.338000000e-07 V_low
+ 8.338010000e-07 V_low
+ 8.339000000e-07 V_low
+ 8.339010000e-07 V_hig
+ 8.340000000e-07 V_hig
+ 8.340010000e-07 V_hig
+ 8.341000000e-07 V_hig
+ 8.341010000e-07 V_hig
+ 8.342000000e-07 V_hig
+ 8.342010000e-07 V_hig
+ 8.343000000e-07 V_hig
+ 8.343010000e-07 V_hig
+ 8.344000000e-07 V_hig
+ 8.344010000e-07 V_hig
+ 8.345000000e-07 V_hig
+ 8.345010000e-07 V_hig
+ 8.346000000e-07 V_hig
+ 8.346010000e-07 V_hig
+ 8.347000000e-07 V_hig
+ 8.347010000e-07 V_hig
+ 8.348000000e-07 V_hig
+ 8.348010000e-07 V_hig
+ 8.349000000e-07 V_hig
+ 8.349010000e-07 V_hig
+ 8.350000000e-07 V_hig
+ 8.350010000e-07 V_hig
+ 8.351000000e-07 V_hig
+ 8.351010000e-07 V_hig
+ 8.352000000e-07 V_hig
+ 8.352010000e-07 V_hig
+ 8.353000000e-07 V_hig
+ 8.353010000e-07 V_hig
+ 8.354000000e-07 V_hig
+ 8.354010000e-07 V_hig
+ 8.355000000e-07 V_hig
+ 8.355010000e-07 V_hig
+ 8.356000000e-07 V_hig
+ 8.356010000e-07 V_hig
+ 8.357000000e-07 V_hig
+ 8.357010000e-07 V_hig
+ 8.358000000e-07 V_hig
+ 8.358010000e-07 V_hig
+ 8.359000000e-07 V_hig
+ 8.359010000e-07 V_low
+ 8.360000000e-07 V_low
+ 8.360010000e-07 V_low
+ 8.361000000e-07 V_low
+ 8.361010000e-07 V_low
+ 8.362000000e-07 V_low
+ 8.362010000e-07 V_low
+ 8.363000000e-07 V_low
+ 8.363010000e-07 V_low
+ 8.364000000e-07 V_low
+ 8.364010000e-07 V_low
+ 8.365000000e-07 V_low
+ 8.365010000e-07 V_low
+ 8.366000000e-07 V_low
+ 8.366010000e-07 V_low
+ 8.367000000e-07 V_low
+ 8.367010000e-07 V_low
+ 8.368000000e-07 V_low
+ 8.368010000e-07 V_low
+ 8.369000000e-07 V_low
+ 8.369010000e-07 V_hig
+ 8.370000000e-07 V_hig
+ 8.370010000e-07 V_hig
+ 8.371000000e-07 V_hig
+ 8.371010000e-07 V_hig
+ 8.372000000e-07 V_hig
+ 8.372010000e-07 V_hig
+ 8.373000000e-07 V_hig
+ 8.373010000e-07 V_hig
+ 8.374000000e-07 V_hig
+ 8.374010000e-07 V_hig
+ 8.375000000e-07 V_hig
+ 8.375010000e-07 V_hig
+ 8.376000000e-07 V_hig
+ 8.376010000e-07 V_hig
+ 8.377000000e-07 V_hig
+ 8.377010000e-07 V_hig
+ 8.378000000e-07 V_hig
+ 8.378010000e-07 V_hig
+ 8.379000000e-07 V_hig
+ 8.379010000e-07 V_low
+ 8.380000000e-07 V_low
+ 8.380010000e-07 V_low
+ 8.381000000e-07 V_low
+ 8.381010000e-07 V_low
+ 8.382000000e-07 V_low
+ 8.382010000e-07 V_low
+ 8.383000000e-07 V_low
+ 8.383010000e-07 V_low
+ 8.384000000e-07 V_low
+ 8.384010000e-07 V_low
+ 8.385000000e-07 V_low
+ 8.385010000e-07 V_low
+ 8.386000000e-07 V_low
+ 8.386010000e-07 V_low
+ 8.387000000e-07 V_low
+ 8.387010000e-07 V_low
+ 8.388000000e-07 V_low
+ 8.388010000e-07 V_low
+ 8.389000000e-07 V_low
+ 8.389010000e-07 V_low
+ 8.390000000e-07 V_low
+ 8.390010000e-07 V_low
+ 8.391000000e-07 V_low
+ 8.391010000e-07 V_low
+ 8.392000000e-07 V_low
+ 8.392010000e-07 V_low
+ 8.393000000e-07 V_low
+ 8.393010000e-07 V_low
+ 8.394000000e-07 V_low
+ 8.394010000e-07 V_low
+ 8.395000000e-07 V_low
+ 8.395010000e-07 V_low
+ 8.396000000e-07 V_low
+ 8.396010000e-07 V_low
+ 8.397000000e-07 V_low
+ 8.397010000e-07 V_low
+ 8.398000000e-07 V_low
+ 8.398010000e-07 V_low
+ 8.399000000e-07 V_low
+ 8.399010000e-07 V_low
+ 8.400000000e-07 V_low
+ 8.400010000e-07 V_low
+ 8.401000000e-07 V_low
+ 8.401010000e-07 V_low
+ 8.402000000e-07 V_low
+ 8.402010000e-07 V_low
+ 8.403000000e-07 V_low
+ 8.403010000e-07 V_low
+ 8.404000000e-07 V_low
+ 8.404010000e-07 V_low
+ 8.405000000e-07 V_low
+ 8.405010000e-07 V_low
+ 8.406000000e-07 V_low
+ 8.406010000e-07 V_low
+ 8.407000000e-07 V_low
+ 8.407010000e-07 V_low
+ 8.408000000e-07 V_low
+ 8.408010000e-07 V_low
+ 8.409000000e-07 V_low
+ 8.409010000e-07 V_hig
+ 8.410000000e-07 V_hig
+ 8.410010000e-07 V_hig
+ 8.411000000e-07 V_hig
+ 8.411010000e-07 V_hig
+ 8.412000000e-07 V_hig
+ 8.412010000e-07 V_hig
+ 8.413000000e-07 V_hig
+ 8.413010000e-07 V_hig
+ 8.414000000e-07 V_hig
+ 8.414010000e-07 V_hig
+ 8.415000000e-07 V_hig
+ 8.415010000e-07 V_hig
+ 8.416000000e-07 V_hig
+ 8.416010000e-07 V_hig
+ 8.417000000e-07 V_hig
+ 8.417010000e-07 V_hig
+ 8.418000000e-07 V_hig
+ 8.418010000e-07 V_hig
+ 8.419000000e-07 V_hig
+ 8.419010000e-07 V_hig
+ 8.420000000e-07 V_hig
+ 8.420010000e-07 V_hig
+ 8.421000000e-07 V_hig
+ 8.421010000e-07 V_hig
+ 8.422000000e-07 V_hig
+ 8.422010000e-07 V_hig
+ 8.423000000e-07 V_hig
+ 8.423010000e-07 V_hig
+ 8.424000000e-07 V_hig
+ 8.424010000e-07 V_hig
+ 8.425000000e-07 V_hig
+ 8.425010000e-07 V_hig
+ 8.426000000e-07 V_hig
+ 8.426010000e-07 V_hig
+ 8.427000000e-07 V_hig
+ 8.427010000e-07 V_hig
+ 8.428000000e-07 V_hig
+ 8.428010000e-07 V_hig
+ 8.429000000e-07 V_hig
+ 8.429010000e-07 V_hig
+ 8.430000000e-07 V_hig
+ 8.430010000e-07 V_hig
+ 8.431000000e-07 V_hig
+ 8.431010000e-07 V_hig
+ 8.432000000e-07 V_hig
+ 8.432010000e-07 V_hig
+ 8.433000000e-07 V_hig
+ 8.433010000e-07 V_hig
+ 8.434000000e-07 V_hig
+ 8.434010000e-07 V_hig
+ 8.435000000e-07 V_hig
+ 8.435010000e-07 V_hig
+ 8.436000000e-07 V_hig
+ 8.436010000e-07 V_hig
+ 8.437000000e-07 V_hig
+ 8.437010000e-07 V_hig
+ 8.438000000e-07 V_hig
+ 8.438010000e-07 V_hig
+ 8.439000000e-07 V_hig
+ 8.439010000e-07 V_hig
+ 8.440000000e-07 V_hig
+ 8.440010000e-07 V_hig
+ 8.441000000e-07 V_hig
+ 8.441010000e-07 V_hig
+ 8.442000000e-07 V_hig
+ 8.442010000e-07 V_hig
+ 8.443000000e-07 V_hig
+ 8.443010000e-07 V_hig
+ 8.444000000e-07 V_hig
+ 8.444010000e-07 V_hig
+ 8.445000000e-07 V_hig
+ 8.445010000e-07 V_hig
+ 8.446000000e-07 V_hig
+ 8.446010000e-07 V_hig
+ 8.447000000e-07 V_hig
+ 8.447010000e-07 V_hig
+ 8.448000000e-07 V_hig
+ 8.448010000e-07 V_hig
+ 8.449000000e-07 V_hig
+ 8.449010000e-07 V_hig
+ 8.450000000e-07 V_hig
+ 8.450010000e-07 V_hig
+ 8.451000000e-07 V_hig
+ 8.451010000e-07 V_hig
+ 8.452000000e-07 V_hig
+ 8.452010000e-07 V_hig
+ 8.453000000e-07 V_hig
+ 8.453010000e-07 V_hig
+ 8.454000000e-07 V_hig
+ 8.454010000e-07 V_hig
+ 8.455000000e-07 V_hig
+ 8.455010000e-07 V_hig
+ 8.456000000e-07 V_hig
+ 8.456010000e-07 V_hig
+ 8.457000000e-07 V_hig
+ 8.457010000e-07 V_hig
+ 8.458000000e-07 V_hig
+ 8.458010000e-07 V_hig
+ 8.459000000e-07 V_hig
+ 8.459010000e-07 V_hig
+ 8.460000000e-07 V_hig
+ 8.460010000e-07 V_hig
+ 8.461000000e-07 V_hig
+ 8.461010000e-07 V_hig
+ 8.462000000e-07 V_hig
+ 8.462010000e-07 V_hig
+ 8.463000000e-07 V_hig
+ 8.463010000e-07 V_hig
+ 8.464000000e-07 V_hig
+ 8.464010000e-07 V_hig
+ 8.465000000e-07 V_hig
+ 8.465010000e-07 V_hig
+ 8.466000000e-07 V_hig
+ 8.466010000e-07 V_hig
+ 8.467000000e-07 V_hig
+ 8.467010000e-07 V_hig
+ 8.468000000e-07 V_hig
+ 8.468010000e-07 V_hig
+ 8.469000000e-07 V_hig
+ 8.469010000e-07 V_hig
+ 8.470000000e-07 V_hig
+ 8.470010000e-07 V_hig
+ 8.471000000e-07 V_hig
+ 8.471010000e-07 V_hig
+ 8.472000000e-07 V_hig
+ 8.472010000e-07 V_hig
+ 8.473000000e-07 V_hig
+ 8.473010000e-07 V_hig
+ 8.474000000e-07 V_hig
+ 8.474010000e-07 V_hig
+ 8.475000000e-07 V_hig
+ 8.475010000e-07 V_hig
+ 8.476000000e-07 V_hig
+ 8.476010000e-07 V_hig
+ 8.477000000e-07 V_hig
+ 8.477010000e-07 V_hig
+ 8.478000000e-07 V_hig
+ 8.478010000e-07 V_hig
+ 8.479000000e-07 V_hig
+ 8.479010000e-07 V_hig
+ 8.480000000e-07 V_hig
+ 8.480010000e-07 V_hig
+ 8.481000000e-07 V_hig
+ 8.481010000e-07 V_hig
+ 8.482000000e-07 V_hig
+ 8.482010000e-07 V_hig
+ 8.483000000e-07 V_hig
+ 8.483010000e-07 V_hig
+ 8.484000000e-07 V_hig
+ 8.484010000e-07 V_hig
+ 8.485000000e-07 V_hig
+ 8.485010000e-07 V_hig
+ 8.486000000e-07 V_hig
+ 8.486010000e-07 V_hig
+ 8.487000000e-07 V_hig
+ 8.487010000e-07 V_hig
+ 8.488000000e-07 V_hig
+ 8.488010000e-07 V_hig
+ 8.489000000e-07 V_hig
+ 8.489010000e-07 V_hig
+ 8.490000000e-07 V_hig
+ 8.490010000e-07 V_hig
+ 8.491000000e-07 V_hig
+ 8.491010000e-07 V_hig
+ 8.492000000e-07 V_hig
+ 8.492010000e-07 V_hig
+ 8.493000000e-07 V_hig
+ 8.493010000e-07 V_hig
+ 8.494000000e-07 V_hig
+ 8.494010000e-07 V_hig
+ 8.495000000e-07 V_hig
+ 8.495010000e-07 V_hig
+ 8.496000000e-07 V_hig
+ 8.496010000e-07 V_hig
+ 8.497000000e-07 V_hig
+ 8.497010000e-07 V_hig
+ 8.498000000e-07 V_hig
+ 8.498010000e-07 V_hig
+ 8.499000000e-07 V_hig
+ 8.499010000e-07 V_low
+ 8.500000000e-07 V_low
+ 8.500010000e-07 V_low
+ 8.501000000e-07 V_low
+ 8.501010000e-07 V_low
+ 8.502000000e-07 V_low
+ 8.502010000e-07 V_low
+ 8.503000000e-07 V_low
+ 8.503010000e-07 V_low
+ 8.504000000e-07 V_low
+ 8.504010000e-07 V_low
+ 8.505000000e-07 V_low
+ 8.505010000e-07 V_low
+ 8.506000000e-07 V_low
+ 8.506010000e-07 V_low
+ 8.507000000e-07 V_low
+ 8.507010000e-07 V_low
+ 8.508000000e-07 V_low
+ 8.508010000e-07 V_low
+ 8.509000000e-07 V_low
+ 8.509010000e-07 V_hig
+ 8.510000000e-07 V_hig
+ 8.510010000e-07 V_hig
+ 8.511000000e-07 V_hig
+ 8.511010000e-07 V_hig
+ 8.512000000e-07 V_hig
+ 8.512010000e-07 V_hig
+ 8.513000000e-07 V_hig
+ 8.513010000e-07 V_hig
+ 8.514000000e-07 V_hig
+ 8.514010000e-07 V_hig
+ 8.515000000e-07 V_hig
+ 8.515010000e-07 V_hig
+ 8.516000000e-07 V_hig
+ 8.516010000e-07 V_hig
+ 8.517000000e-07 V_hig
+ 8.517010000e-07 V_hig
+ 8.518000000e-07 V_hig
+ 8.518010000e-07 V_hig
+ 8.519000000e-07 V_hig
+ 8.519010000e-07 V_hig
+ 8.520000000e-07 V_hig
+ 8.520010000e-07 V_hig
+ 8.521000000e-07 V_hig
+ 8.521010000e-07 V_hig
+ 8.522000000e-07 V_hig
+ 8.522010000e-07 V_hig
+ 8.523000000e-07 V_hig
+ 8.523010000e-07 V_hig
+ 8.524000000e-07 V_hig
+ 8.524010000e-07 V_hig
+ 8.525000000e-07 V_hig
+ 8.525010000e-07 V_hig
+ 8.526000000e-07 V_hig
+ 8.526010000e-07 V_hig
+ 8.527000000e-07 V_hig
+ 8.527010000e-07 V_hig
+ 8.528000000e-07 V_hig
+ 8.528010000e-07 V_hig
+ 8.529000000e-07 V_hig
+ 8.529010000e-07 V_hig
+ 8.530000000e-07 V_hig
+ 8.530010000e-07 V_hig
+ 8.531000000e-07 V_hig
+ 8.531010000e-07 V_hig
+ 8.532000000e-07 V_hig
+ 8.532010000e-07 V_hig
+ 8.533000000e-07 V_hig
+ 8.533010000e-07 V_hig
+ 8.534000000e-07 V_hig
+ 8.534010000e-07 V_hig
+ 8.535000000e-07 V_hig
+ 8.535010000e-07 V_hig
+ 8.536000000e-07 V_hig
+ 8.536010000e-07 V_hig
+ 8.537000000e-07 V_hig
+ 8.537010000e-07 V_hig
+ 8.538000000e-07 V_hig
+ 8.538010000e-07 V_hig
+ 8.539000000e-07 V_hig
+ 8.539010000e-07 V_low
+ 8.540000000e-07 V_low
+ 8.540010000e-07 V_low
+ 8.541000000e-07 V_low
+ 8.541010000e-07 V_low
+ 8.542000000e-07 V_low
+ 8.542010000e-07 V_low
+ 8.543000000e-07 V_low
+ 8.543010000e-07 V_low
+ 8.544000000e-07 V_low
+ 8.544010000e-07 V_low
+ 8.545000000e-07 V_low
+ 8.545010000e-07 V_low
+ 8.546000000e-07 V_low
+ 8.546010000e-07 V_low
+ 8.547000000e-07 V_low
+ 8.547010000e-07 V_low
+ 8.548000000e-07 V_low
+ 8.548010000e-07 V_low
+ 8.549000000e-07 V_low
+ 8.549010000e-07 V_hig
+ 8.550000000e-07 V_hig
+ 8.550010000e-07 V_hig
+ 8.551000000e-07 V_hig
+ 8.551010000e-07 V_hig
+ 8.552000000e-07 V_hig
+ 8.552010000e-07 V_hig
+ 8.553000000e-07 V_hig
+ 8.553010000e-07 V_hig
+ 8.554000000e-07 V_hig
+ 8.554010000e-07 V_hig
+ 8.555000000e-07 V_hig
+ 8.555010000e-07 V_hig
+ 8.556000000e-07 V_hig
+ 8.556010000e-07 V_hig
+ 8.557000000e-07 V_hig
+ 8.557010000e-07 V_hig
+ 8.558000000e-07 V_hig
+ 8.558010000e-07 V_hig
+ 8.559000000e-07 V_hig
+ 8.559010000e-07 V_hig
+ 8.560000000e-07 V_hig
+ 8.560010000e-07 V_hig
+ 8.561000000e-07 V_hig
+ 8.561010000e-07 V_hig
+ 8.562000000e-07 V_hig
+ 8.562010000e-07 V_hig
+ 8.563000000e-07 V_hig
+ 8.563010000e-07 V_hig
+ 8.564000000e-07 V_hig
+ 8.564010000e-07 V_hig
+ 8.565000000e-07 V_hig
+ 8.565010000e-07 V_hig
+ 8.566000000e-07 V_hig
+ 8.566010000e-07 V_hig
+ 8.567000000e-07 V_hig
+ 8.567010000e-07 V_hig
+ 8.568000000e-07 V_hig
+ 8.568010000e-07 V_hig
+ 8.569000000e-07 V_hig
+ 8.569010000e-07 V_low
+ 8.570000000e-07 V_low
+ 8.570010000e-07 V_low
+ 8.571000000e-07 V_low
+ 8.571010000e-07 V_low
+ 8.572000000e-07 V_low
+ 8.572010000e-07 V_low
+ 8.573000000e-07 V_low
+ 8.573010000e-07 V_low
+ 8.574000000e-07 V_low
+ 8.574010000e-07 V_low
+ 8.575000000e-07 V_low
+ 8.575010000e-07 V_low
+ 8.576000000e-07 V_low
+ 8.576010000e-07 V_low
+ 8.577000000e-07 V_low
+ 8.577010000e-07 V_low
+ 8.578000000e-07 V_low
+ 8.578010000e-07 V_low
+ 8.579000000e-07 V_low
+ 8.579010000e-07 V_low
+ 8.580000000e-07 V_low
+ 8.580010000e-07 V_low
+ 8.581000000e-07 V_low
+ 8.581010000e-07 V_low
+ 8.582000000e-07 V_low
+ 8.582010000e-07 V_low
+ 8.583000000e-07 V_low
+ 8.583010000e-07 V_low
+ 8.584000000e-07 V_low
+ 8.584010000e-07 V_low
+ 8.585000000e-07 V_low
+ 8.585010000e-07 V_low
+ 8.586000000e-07 V_low
+ 8.586010000e-07 V_low
+ 8.587000000e-07 V_low
+ 8.587010000e-07 V_low
+ 8.588000000e-07 V_low
+ 8.588010000e-07 V_low
+ 8.589000000e-07 V_low
+ 8.589010000e-07 V_low
+ 8.590000000e-07 V_low
+ 8.590010000e-07 V_low
+ 8.591000000e-07 V_low
+ 8.591010000e-07 V_low
+ 8.592000000e-07 V_low
+ 8.592010000e-07 V_low
+ 8.593000000e-07 V_low
+ 8.593010000e-07 V_low
+ 8.594000000e-07 V_low
+ 8.594010000e-07 V_low
+ 8.595000000e-07 V_low
+ 8.595010000e-07 V_low
+ 8.596000000e-07 V_low
+ 8.596010000e-07 V_low
+ 8.597000000e-07 V_low
+ 8.597010000e-07 V_low
+ 8.598000000e-07 V_low
+ 8.598010000e-07 V_low
+ 8.599000000e-07 V_low
+ 8.599010000e-07 V_hig
+ 8.600000000e-07 V_hig
+ 8.600010000e-07 V_hig
+ 8.601000000e-07 V_hig
+ 8.601010000e-07 V_hig
+ 8.602000000e-07 V_hig
+ 8.602010000e-07 V_hig
+ 8.603000000e-07 V_hig
+ 8.603010000e-07 V_hig
+ 8.604000000e-07 V_hig
+ 8.604010000e-07 V_hig
+ 8.605000000e-07 V_hig
+ 8.605010000e-07 V_hig
+ 8.606000000e-07 V_hig
+ 8.606010000e-07 V_hig
+ 8.607000000e-07 V_hig
+ 8.607010000e-07 V_hig
+ 8.608000000e-07 V_hig
+ 8.608010000e-07 V_hig
+ 8.609000000e-07 V_hig
+ 8.609010000e-07 V_hig
+ 8.610000000e-07 V_hig
+ 8.610010000e-07 V_hig
+ 8.611000000e-07 V_hig
+ 8.611010000e-07 V_hig
+ 8.612000000e-07 V_hig
+ 8.612010000e-07 V_hig
+ 8.613000000e-07 V_hig
+ 8.613010000e-07 V_hig
+ 8.614000000e-07 V_hig
+ 8.614010000e-07 V_hig
+ 8.615000000e-07 V_hig
+ 8.615010000e-07 V_hig
+ 8.616000000e-07 V_hig
+ 8.616010000e-07 V_hig
+ 8.617000000e-07 V_hig
+ 8.617010000e-07 V_hig
+ 8.618000000e-07 V_hig
+ 8.618010000e-07 V_hig
+ 8.619000000e-07 V_hig
+ 8.619010000e-07 V_low
+ 8.620000000e-07 V_low
+ 8.620010000e-07 V_low
+ 8.621000000e-07 V_low
+ 8.621010000e-07 V_low
+ 8.622000000e-07 V_low
+ 8.622010000e-07 V_low
+ 8.623000000e-07 V_low
+ 8.623010000e-07 V_low
+ 8.624000000e-07 V_low
+ 8.624010000e-07 V_low
+ 8.625000000e-07 V_low
+ 8.625010000e-07 V_low
+ 8.626000000e-07 V_low
+ 8.626010000e-07 V_low
+ 8.627000000e-07 V_low
+ 8.627010000e-07 V_low
+ 8.628000000e-07 V_low
+ 8.628010000e-07 V_low
+ 8.629000000e-07 V_low
+ 8.629010000e-07 V_low
+ 8.630000000e-07 V_low
+ 8.630010000e-07 V_low
+ 8.631000000e-07 V_low
+ 8.631010000e-07 V_low
+ 8.632000000e-07 V_low
+ 8.632010000e-07 V_low
+ 8.633000000e-07 V_low
+ 8.633010000e-07 V_low
+ 8.634000000e-07 V_low
+ 8.634010000e-07 V_low
+ 8.635000000e-07 V_low
+ 8.635010000e-07 V_low
+ 8.636000000e-07 V_low
+ 8.636010000e-07 V_low
+ 8.637000000e-07 V_low
+ 8.637010000e-07 V_low
+ 8.638000000e-07 V_low
+ 8.638010000e-07 V_low
+ 8.639000000e-07 V_low
+ 8.639010000e-07 V_low
+ 8.640000000e-07 V_low
+ 8.640010000e-07 V_low
+ 8.641000000e-07 V_low
+ 8.641010000e-07 V_low
+ 8.642000000e-07 V_low
+ 8.642010000e-07 V_low
+ 8.643000000e-07 V_low
+ 8.643010000e-07 V_low
+ 8.644000000e-07 V_low
+ 8.644010000e-07 V_low
+ 8.645000000e-07 V_low
+ 8.645010000e-07 V_low
+ 8.646000000e-07 V_low
+ 8.646010000e-07 V_low
+ 8.647000000e-07 V_low
+ 8.647010000e-07 V_low
+ 8.648000000e-07 V_low
+ 8.648010000e-07 V_low
+ 8.649000000e-07 V_low
+ 8.649010000e-07 V_low
+ 8.650000000e-07 V_low
+ 8.650010000e-07 V_low
+ 8.651000000e-07 V_low
+ 8.651010000e-07 V_low
+ 8.652000000e-07 V_low
+ 8.652010000e-07 V_low
+ 8.653000000e-07 V_low
+ 8.653010000e-07 V_low
+ 8.654000000e-07 V_low
+ 8.654010000e-07 V_low
+ 8.655000000e-07 V_low
+ 8.655010000e-07 V_low
+ 8.656000000e-07 V_low
+ 8.656010000e-07 V_low
+ 8.657000000e-07 V_low
+ 8.657010000e-07 V_low
+ 8.658000000e-07 V_low
+ 8.658010000e-07 V_low
+ 8.659000000e-07 V_low
+ 8.659010000e-07 V_hig
+ 8.660000000e-07 V_hig
+ 8.660010000e-07 V_hig
+ 8.661000000e-07 V_hig
+ 8.661010000e-07 V_hig
+ 8.662000000e-07 V_hig
+ 8.662010000e-07 V_hig
+ 8.663000000e-07 V_hig
+ 8.663010000e-07 V_hig
+ 8.664000000e-07 V_hig
+ 8.664010000e-07 V_hig
+ 8.665000000e-07 V_hig
+ 8.665010000e-07 V_hig
+ 8.666000000e-07 V_hig
+ 8.666010000e-07 V_hig
+ 8.667000000e-07 V_hig
+ 8.667010000e-07 V_hig
+ 8.668000000e-07 V_hig
+ 8.668010000e-07 V_hig
+ 8.669000000e-07 V_hig
+ 8.669010000e-07 V_low
+ 8.670000000e-07 V_low
+ 8.670010000e-07 V_low
+ 8.671000000e-07 V_low
+ 8.671010000e-07 V_low
+ 8.672000000e-07 V_low
+ 8.672010000e-07 V_low
+ 8.673000000e-07 V_low
+ 8.673010000e-07 V_low
+ 8.674000000e-07 V_low
+ 8.674010000e-07 V_low
+ 8.675000000e-07 V_low
+ 8.675010000e-07 V_low
+ 8.676000000e-07 V_low
+ 8.676010000e-07 V_low
+ 8.677000000e-07 V_low
+ 8.677010000e-07 V_low
+ 8.678000000e-07 V_low
+ 8.678010000e-07 V_low
+ 8.679000000e-07 V_low
+ 8.679010000e-07 V_hig
+ 8.680000000e-07 V_hig
+ 8.680010000e-07 V_hig
+ 8.681000000e-07 V_hig
+ 8.681010000e-07 V_hig
+ 8.682000000e-07 V_hig
+ 8.682010000e-07 V_hig
+ 8.683000000e-07 V_hig
+ 8.683010000e-07 V_hig
+ 8.684000000e-07 V_hig
+ 8.684010000e-07 V_hig
+ 8.685000000e-07 V_hig
+ 8.685010000e-07 V_hig
+ 8.686000000e-07 V_hig
+ 8.686010000e-07 V_hig
+ 8.687000000e-07 V_hig
+ 8.687010000e-07 V_hig
+ 8.688000000e-07 V_hig
+ 8.688010000e-07 V_hig
+ 8.689000000e-07 V_hig
+ 8.689010000e-07 V_low
+ 8.690000000e-07 V_low
+ 8.690010000e-07 V_low
+ 8.691000000e-07 V_low
+ 8.691010000e-07 V_low
+ 8.692000000e-07 V_low
+ 8.692010000e-07 V_low
+ 8.693000000e-07 V_low
+ 8.693010000e-07 V_low
+ 8.694000000e-07 V_low
+ 8.694010000e-07 V_low
+ 8.695000000e-07 V_low
+ 8.695010000e-07 V_low
+ 8.696000000e-07 V_low
+ 8.696010000e-07 V_low
+ 8.697000000e-07 V_low
+ 8.697010000e-07 V_low
+ 8.698000000e-07 V_low
+ 8.698010000e-07 V_low
+ 8.699000000e-07 V_low
+ 8.699010000e-07 V_hig
+ 8.700000000e-07 V_hig
+ 8.700010000e-07 V_hig
+ 8.701000000e-07 V_hig
+ 8.701010000e-07 V_hig
+ 8.702000000e-07 V_hig
+ 8.702010000e-07 V_hig
+ 8.703000000e-07 V_hig
+ 8.703010000e-07 V_hig
+ 8.704000000e-07 V_hig
+ 8.704010000e-07 V_hig
+ 8.705000000e-07 V_hig
+ 8.705010000e-07 V_hig
+ 8.706000000e-07 V_hig
+ 8.706010000e-07 V_hig
+ 8.707000000e-07 V_hig
+ 8.707010000e-07 V_hig
+ 8.708000000e-07 V_hig
+ 8.708010000e-07 V_hig
+ 8.709000000e-07 V_hig
+ 8.709010000e-07 V_hig
+ 8.710000000e-07 V_hig
+ 8.710010000e-07 V_hig
+ 8.711000000e-07 V_hig
+ 8.711010000e-07 V_hig
+ 8.712000000e-07 V_hig
+ 8.712010000e-07 V_hig
+ 8.713000000e-07 V_hig
+ 8.713010000e-07 V_hig
+ 8.714000000e-07 V_hig
+ 8.714010000e-07 V_hig
+ 8.715000000e-07 V_hig
+ 8.715010000e-07 V_hig
+ 8.716000000e-07 V_hig
+ 8.716010000e-07 V_hig
+ 8.717000000e-07 V_hig
+ 8.717010000e-07 V_hig
+ 8.718000000e-07 V_hig
+ 8.718010000e-07 V_hig
+ 8.719000000e-07 V_hig
+ 8.719010000e-07 V_hig
+ 8.720000000e-07 V_hig
+ 8.720010000e-07 V_hig
+ 8.721000000e-07 V_hig
+ 8.721010000e-07 V_hig
+ 8.722000000e-07 V_hig
+ 8.722010000e-07 V_hig
+ 8.723000000e-07 V_hig
+ 8.723010000e-07 V_hig
+ 8.724000000e-07 V_hig
+ 8.724010000e-07 V_hig
+ 8.725000000e-07 V_hig
+ 8.725010000e-07 V_hig
+ 8.726000000e-07 V_hig
+ 8.726010000e-07 V_hig
+ 8.727000000e-07 V_hig
+ 8.727010000e-07 V_hig
+ 8.728000000e-07 V_hig
+ 8.728010000e-07 V_hig
+ 8.729000000e-07 V_hig
+ 8.729010000e-07 V_hig
+ 8.730000000e-07 V_hig
+ 8.730010000e-07 V_hig
+ 8.731000000e-07 V_hig
+ 8.731010000e-07 V_hig
+ 8.732000000e-07 V_hig
+ 8.732010000e-07 V_hig
+ 8.733000000e-07 V_hig
+ 8.733010000e-07 V_hig
+ 8.734000000e-07 V_hig
+ 8.734010000e-07 V_hig
+ 8.735000000e-07 V_hig
+ 8.735010000e-07 V_hig
+ 8.736000000e-07 V_hig
+ 8.736010000e-07 V_hig
+ 8.737000000e-07 V_hig
+ 8.737010000e-07 V_hig
+ 8.738000000e-07 V_hig
+ 8.738010000e-07 V_hig
+ 8.739000000e-07 V_hig
+ 8.739010000e-07 V_hig
+ 8.740000000e-07 V_hig
+ 8.740010000e-07 V_hig
+ 8.741000000e-07 V_hig
+ 8.741010000e-07 V_hig
+ 8.742000000e-07 V_hig
+ 8.742010000e-07 V_hig
+ 8.743000000e-07 V_hig
+ 8.743010000e-07 V_hig
+ 8.744000000e-07 V_hig
+ 8.744010000e-07 V_hig
+ 8.745000000e-07 V_hig
+ 8.745010000e-07 V_hig
+ 8.746000000e-07 V_hig
+ 8.746010000e-07 V_hig
+ 8.747000000e-07 V_hig
+ 8.747010000e-07 V_hig
+ 8.748000000e-07 V_hig
+ 8.748010000e-07 V_hig
+ 8.749000000e-07 V_hig
+ 8.749010000e-07 V_hig
+ 8.750000000e-07 V_hig
+ 8.750010000e-07 V_hig
+ 8.751000000e-07 V_hig
+ 8.751010000e-07 V_hig
+ 8.752000000e-07 V_hig
+ 8.752010000e-07 V_hig
+ 8.753000000e-07 V_hig
+ 8.753010000e-07 V_hig
+ 8.754000000e-07 V_hig
+ 8.754010000e-07 V_hig
+ 8.755000000e-07 V_hig
+ 8.755010000e-07 V_hig
+ 8.756000000e-07 V_hig
+ 8.756010000e-07 V_hig
+ 8.757000000e-07 V_hig
+ 8.757010000e-07 V_hig
+ 8.758000000e-07 V_hig
+ 8.758010000e-07 V_hig
+ 8.759000000e-07 V_hig
+ 8.759010000e-07 V_low
+ 8.760000000e-07 V_low
+ 8.760010000e-07 V_low
+ 8.761000000e-07 V_low
+ 8.761010000e-07 V_low
+ 8.762000000e-07 V_low
+ 8.762010000e-07 V_low
+ 8.763000000e-07 V_low
+ 8.763010000e-07 V_low
+ 8.764000000e-07 V_low
+ 8.764010000e-07 V_low
+ 8.765000000e-07 V_low
+ 8.765010000e-07 V_low
+ 8.766000000e-07 V_low
+ 8.766010000e-07 V_low
+ 8.767000000e-07 V_low
+ 8.767010000e-07 V_low
+ 8.768000000e-07 V_low
+ 8.768010000e-07 V_low
+ 8.769000000e-07 V_low
+ 8.769010000e-07 V_low
+ 8.770000000e-07 V_low
+ 8.770010000e-07 V_low
+ 8.771000000e-07 V_low
+ 8.771010000e-07 V_low
+ 8.772000000e-07 V_low
+ 8.772010000e-07 V_low
+ 8.773000000e-07 V_low
+ 8.773010000e-07 V_low
+ 8.774000000e-07 V_low
+ 8.774010000e-07 V_low
+ 8.775000000e-07 V_low
+ 8.775010000e-07 V_low
+ 8.776000000e-07 V_low
+ 8.776010000e-07 V_low
+ 8.777000000e-07 V_low
+ 8.777010000e-07 V_low
+ 8.778000000e-07 V_low
+ 8.778010000e-07 V_low
+ 8.779000000e-07 V_low
+ 8.779010000e-07 V_hig
+ 8.780000000e-07 V_hig
+ 8.780010000e-07 V_hig
+ 8.781000000e-07 V_hig
+ 8.781010000e-07 V_hig
+ 8.782000000e-07 V_hig
+ 8.782010000e-07 V_hig
+ 8.783000000e-07 V_hig
+ 8.783010000e-07 V_hig
+ 8.784000000e-07 V_hig
+ 8.784010000e-07 V_hig
+ 8.785000000e-07 V_hig
+ 8.785010000e-07 V_hig
+ 8.786000000e-07 V_hig
+ 8.786010000e-07 V_hig
+ 8.787000000e-07 V_hig
+ 8.787010000e-07 V_hig
+ 8.788000000e-07 V_hig
+ 8.788010000e-07 V_hig
+ 8.789000000e-07 V_hig
+ 8.789010000e-07 V_hig
+ 8.790000000e-07 V_hig
+ 8.790010000e-07 V_hig
+ 8.791000000e-07 V_hig
+ 8.791010000e-07 V_hig
+ 8.792000000e-07 V_hig
+ 8.792010000e-07 V_hig
+ 8.793000000e-07 V_hig
+ 8.793010000e-07 V_hig
+ 8.794000000e-07 V_hig
+ 8.794010000e-07 V_hig
+ 8.795000000e-07 V_hig
+ 8.795010000e-07 V_hig
+ 8.796000000e-07 V_hig
+ 8.796010000e-07 V_hig
+ 8.797000000e-07 V_hig
+ 8.797010000e-07 V_hig
+ 8.798000000e-07 V_hig
+ 8.798010000e-07 V_hig
+ 8.799000000e-07 V_hig
+ 8.799010000e-07 V_low
+ 8.800000000e-07 V_low
+ 8.800010000e-07 V_low
+ 8.801000000e-07 V_low
+ 8.801010000e-07 V_low
+ 8.802000000e-07 V_low
+ 8.802010000e-07 V_low
+ 8.803000000e-07 V_low
+ 8.803010000e-07 V_low
+ 8.804000000e-07 V_low
+ 8.804010000e-07 V_low
+ 8.805000000e-07 V_low
+ 8.805010000e-07 V_low
+ 8.806000000e-07 V_low
+ 8.806010000e-07 V_low
+ 8.807000000e-07 V_low
+ 8.807010000e-07 V_low
+ 8.808000000e-07 V_low
+ 8.808010000e-07 V_low
+ 8.809000000e-07 V_low
+ 8.809010000e-07 V_low
+ 8.810000000e-07 V_low
+ 8.810010000e-07 V_low
+ 8.811000000e-07 V_low
+ 8.811010000e-07 V_low
+ 8.812000000e-07 V_low
+ 8.812010000e-07 V_low
+ 8.813000000e-07 V_low
+ 8.813010000e-07 V_low
+ 8.814000000e-07 V_low
+ 8.814010000e-07 V_low
+ 8.815000000e-07 V_low
+ 8.815010000e-07 V_low
+ 8.816000000e-07 V_low
+ 8.816010000e-07 V_low
+ 8.817000000e-07 V_low
+ 8.817010000e-07 V_low
+ 8.818000000e-07 V_low
+ 8.818010000e-07 V_low
+ 8.819000000e-07 V_low
+ 8.819010000e-07 V_low
+ 8.820000000e-07 V_low
+ 8.820010000e-07 V_low
+ 8.821000000e-07 V_low
+ 8.821010000e-07 V_low
+ 8.822000000e-07 V_low
+ 8.822010000e-07 V_low
+ 8.823000000e-07 V_low
+ 8.823010000e-07 V_low
+ 8.824000000e-07 V_low
+ 8.824010000e-07 V_low
+ 8.825000000e-07 V_low
+ 8.825010000e-07 V_low
+ 8.826000000e-07 V_low
+ 8.826010000e-07 V_low
+ 8.827000000e-07 V_low
+ 8.827010000e-07 V_low
+ 8.828000000e-07 V_low
+ 8.828010000e-07 V_low
+ 8.829000000e-07 V_low
+ 8.829010000e-07 V_hig
+ 8.830000000e-07 V_hig
+ 8.830010000e-07 V_hig
+ 8.831000000e-07 V_hig
+ 8.831010000e-07 V_hig
+ 8.832000000e-07 V_hig
+ 8.832010000e-07 V_hig
+ 8.833000000e-07 V_hig
+ 8.833010000e-07 V_hig
+ 8.834000000e-07 V_hig
+ 8.834010000e-07 V_hig
+ 8.835000000e-07 V_hig
+ 8.835010000e-07 V_hig
+ 8.836000000e-07 V_hig
+ 8.836010000e-07 V_hig
+ 8.837000000e-07 V_hig
+ 8.837010000e-07 V_hig
+ 8.838000000e-07 V_hig
+ 8.838010000e-07 V_hig
+ 8.839000000e-07 V_hig
+ 8.839010000e-07 V_low
+ 8.840000000e-07 V_low
+ 8.840010000e-07 V_low
+ 8.841000000e-07 V_low
+ 8.841010000e-07 V_low
+ 8.842000000e-07 V_low
+ 8.842010000e-07 V_low
+ 8.843000000e-07 V_low
+ 8.843010000e-07 V_low
+ 8.844000000e-07 V_low
+ 8.844010000e-07 V_low
+ 8.845000000e-07 V_low
+ 8.845010000e-07 V_low
+ 8.846000000e-07 V_low
+ 8.846010000e-07 V_low
+ 8.847000000e-07 V_low
+ 8.847010000e-07 V_low
+ 8.848000000e-07 V_low
+ 8.848010000e-07 V_low
+ 8.849000000e-07 V_low
+ 8.849010000e-07 V_hig
+ 8.850000000e-07 V_hig
+ 8.850010000e-07 V_hig
+ 8.851000000e-07 V_hig
+ 8.851010000e-07 V_hig
+ 8.852000000e-07 V_hig
+ 8.852010000e-07 V_hig
+ 8.853000000e-07 V_hig
+ 8.853010000e-07 V_hig
+ 8.854000000e-07 V_hig
+ 8.854010000e-07 V_hig
+ 8.855000000e-07 V_hig
+ 8.855010000e-07 V_hig
+ 8.856000000e-07 V_hig
+ 8.856010000e-07 V_hig
+ 8.857000000e-07 V_hig
+ 8.857010000e-07 V_hig
+ 8.858000000e-07 V_hig
+ 8.858010000e-07 V_hig
+ 8.859000000e-07 V_hig
+ 8.859010000e-07 V_low
+ 8.860000000e-07 V_low
+ 8.860010000e-07 V_low
+ 8.861000000e-07 V_low
+ 8.861010000e-07 V_low
+ 8.862000000e-07 V_low
+ 8.862010000e-07 V_low
+ 8.863000000e-07 V_low
+ 8.863010000e-07 V_low
+ 8.864000000e-07 V_low
+ 8.864010000e-07 V_low
+ 8.865000000e-07 V_low
+ 8.865010000e-07 V_low
+ 8.866000000e-07 V_low
+ 8.866010000e-07 V_low
+ 8.867000000e-07 V_low
+ 8.867010000e-07 V_low
+ 8.868000000e-07 V_low
+ 8.868010000e-07 V_low
+ 8.869000000e-07 V_low
+ 8.869010000e-07 V_low
+ 8.870000000e-07 V_low
+ 8.870010000e-07 V_low
+ 8.871000000e-07 V_low
+ 8.871010000e-07 V_low
+ 8.872000000e-07 V_low
+ 8.872010000e-07 V_low
+ 8.873000000e-07 V_low
+ 8.873010000e-07 V_low
+ 8.874000000e-07 V_low
+ 8.874010000e-07 V_low
+ 8.875000000e-07 V_low
+ 8.875010000e-07 V_low
+ 8.876000000e-07 V_low
+ 8.876010000e-07 V_low
+ 8.877000000e-07 V_low
+ 8.877010000e-07 V_low
+ 8.878000000e-07 V_low
+ 8.878010000e-07 V_low
+ 8.879000000e-07 V_low
+ 8.879010000e-07 V_hig
+ 8.880000000e-07 V_hig
+ 8.880010000e-07 V_hig
+ 8.881000000e-07 V_hig
+ 8.881010000e-07 V_hig
+ 8.882000000e-07 V_hig
+ 8.882010000e-07 V_hig
+ 8.883000000e-07 V_hig
+ 8.883010000e-07 V_hig
+ 8.884000000e-07 V_hig
+ 8.884010000e-07 V_hig
+ 8.885000000e-07 V_hig
+ 8.885010000e-07 V_hig
+ 8.886000000e-07 V_hig
+ 8.886010000e-07 V_hig
+ 8.887000000e-07 V_hig
+ 8.887010000e-07 V_hig
+ 8.888000000e-07 V_hig
+ 8.888010000e-07 V_hig
+ 8.889000000e-07 V_hig
+ 8.889010000e-07 V_hig
+ 8.890000000e-07 V_hig
+ 8.890010000e-07 V_hig
+ 8.891000000e-07 V_hig
+ 8.891010000e-07 V_hig
+ 8.892000000e-07 V_hig
+ 8.892010000e-07 V_hig
+ 8.893000000e-07 V_hig
+ 8.893010000e-07 V_hig
+ 8.894000000e-07 V_hig
+ 8.894010000e-07 V_hig
+ 8.895000000e-07 V_hig
+ 8.895010000e-07 V_hig
+ 8.896000000e-07 V_hig
+ 8.896010000e-07 V_hig
+ 8.897000000e-07 V_hig
+ 8.897010000e-07 V_hig
+ 8.898000000e-07 V_hig
+ 8.898010000e-07 V_hig
+ 8.899000000e-07 V_hig
+ 8.899010000e-07 V_hig
+ 8.900000000e-07 V_hig
+ 8.900010000e-07 V_hig
+ 8.901000000e-07 V_hig
+ 8.901010000e-07 V_hig
+ 8.902000000e-07 V_hig
+ 8.902010000e-07 V_hig
+ 8.903000000e-07 V_hig
+ 8.903010000e-07 V_hig
+ 8.904000000e-07 V_hig
+ 8.904010000e-07 V_hig
+ 8.905000000e-07 V_hig
+ 8.905010000e-07 V_hig
+ 8.906000000e-07 V_hig
+ 8.906010000e-07 V_hig
+ 8.907000000e-07 V_hig
+ 8.907010000e-07 V_hig
+ 8.908000000e-07 V_hig
+ 8.908010000e-07 V_hig
+ 8.909000000e-07 V_hig
+ 8.909010000e-07 V_hig
+ 8.910000000e-07 V_hig
+ 8.910010000e-07 V_hig
+ 8.911000000e-07 V_hig
+ 8.911010000e-07 V_hig
+ 8.912000000e-07 V_hig
+ 8.912010000e-07 V_hig
+ 8.913000000e-07 V_hig
+ 8.913010000e-07 V_hig
+ 8.914000000e-07 V_hig
+ 8.914010000e-07 V_hig
+ 8.915000000e-07 V_hig
+ 8.915010000e-07 V_hig
+ 8.916000000e-07 V_hig
+ 8.916010000e-07 V_hig
+ 8.917000000e-07 V_hig
+ 8.917010000e-07 V_hig
+ 8.918000000e-07 V_hig
+ 8.918010000e-07 V_hig
+ 8.919000000e-07 V_hig
+ 8.919010000e-07 V_low
+ 8.920000000e-07 V_low
+ 8.920010000e-07 V_low
+ 8.921000000e-07 V_low
+ 8.921010000e-07 V_low
+ 8.922000000e-07 V_low
+ 8.922010000e-07 V_low
+ 8.923000000e-07 V_low
+ 8.923010000e-07 V_low
+ 8.924000000e-07 V_low
+ 8.924010000e-07 V_low
+ 8.925000000e-07 V_low
+ 8.925010000e-07 V_low
+ 8.926000000e-07 V_low
+ 8.926010000e-07 V_low
+ 8.927000000e-07 V_low
+ 8.927010000e-07 V_low
+ 8.928000000e-07 V_low
+ 8.928010000e-07 V_low
+ 8.929000000e-07 V_low
+ 8.929010000e-07 V_hig
+ 8.930000000e-07 V_hig
+ 8.930010000e-07 V_hig
+ 8.931000000e-07 V_hig
+ 8.931010000e-07 V_hig
+ 8.932000000e-07 V_hig
+ 8.932010000e-07 V_hig
+ 8.933000000e-07 V_hig
+ 8.933010000e-07 V_hig
+ 8.934000000e-07 V_hig
+ 8.934010000e-07 V_hig
+ 8.935000000e-07 V_hig
+ 8.935010000e-07 V_hig
+ 8.936000000e-07 V_hig
+ 8.936010000e-07 V_hig
+ 8.937000000e-07 V_hig
+ 8.937010000e-07 V_hig
+ 8.938000000e-07 V_hig
+ 8.938010000e-07 V_hig
+ 8.939000000e-07 V_hig
+ 8.939010000e-07 V_hig
+ 8.940000000e-07 V_hig
+ 8.940010000e-07 V_hig
+ 8.941000000e-07 V_hig
+ 8.941010000e-07 V_hig
+ 8.942000000e-07 V_hig
+ 8.942010000e-07 V_hig
+ 8.943000000e-07 V_hig
+ 8.943010000e-07 V_hig
+ 8.944000000e-07 V_hig
+ 8.944010000e-07 V_hig
+ 8.945000000e-07 V_hig
+ 8.945010000e-07 V_hig
+ 8.946000000e-07 V_hig
+ 8.946010000e-07 V_hig
+ 8.947000000e-07 V_hig
+ 8.947010000e-07 V_hig
+ 8.948000000e-07 V_hig
+ 8.948010000e-07 V_hig
+ 8.949000000e-07 V_hig
+ 8.949010000e-07 V_low
+ 8.950000000e-07 V_low
+ 8.950010000e-07 V_low
+ 8.951000000e-07 V_low
+ 8.951010000e-07 V_low
+ 8.952000000e-07 V_low
+ 8.952010000e-07 V_low
+ 8.953000000e-07 V_low
+ 8.953010000e-07 V_low
+ 8.954000000e-07 V_low
+ 8.954010000e-07 V_low
+ 8.955000000e-07 V_low
+ 8.955010000e-07 V_low
+ 8.956000000e-07 V_low
+ 8.956010000e-07 V_low
+ 8.957000000e-07 V_low
+ 8.957010000e-07 V_low
+ 8.958000000e-07 V_low
+ 8.958010000e-07 V_low
+ 8.959000000e-07 V_low
+ 8.959010000e-07 V_hig
+ 8.960000000e-07 V_hig
+ 8.960010000e-07 V_hig
+ 8.961000000e-07 V_hig
+ 8.961010000e-07 V_hig
+ 8.962000000e-07 V_hig
+ 8.962010000e-07 V_hig
+ 8.963000000e-07 V_hig
+ 8.963010000e-07 V_hig
+ 8.964000000e-07 V_hig
+ 8.964010000e-07 V_hig
+ 8.965000000e-07 V_hig
+ 8.965010000e-07 V_hig
+ 8.966000000e-07 V_hig
+ 8.966010000e-07 V_hig
+ 8.967000000e-07 V_hig
+ 8.967010000e-07 V_hig
+ 8.968000000e-07 V_hig
+ 8.968010000e-07 V_hig
+ 8.969000000e-07 V_hig
+ 8.969010000e-07 V_hig
+ 8.970000000e-07 V_hig
+ 8.970010000e-07 V_hig
+ 8.971000000e-07 V_hig
+ 8.971010000e-07 V_hig
+ 8.972000000e-07 V_hig
+ 8.972010000e-07 V_hig
+ 8.973000000e-07 V_hig
+ 8.973010000e-07 V_hig
+ 8.974000000e-07 V_hig
+ 8.974010000e-07 V_hig
+ 8.975000000e-07 V_hig
+ 8.975010000e-07 V_hig
+ 8.976000000e-07 V_hig
+ 8.976010000e-07 V_hig
+ 8.977000000e-07 V_hig
+ 8.977010000e-07 V_hig
+ 8.978000000e-07 V_hig
+ 8.978010000e-07 V_hig
+ 8.979000000e-07 V_hig
+ 8.979010000e-07 V_low
+ 8.980000000e-07 V_low
+ 8.980010000e-07 V_low
+ 8.981000000e-07 V_low
+ 8.981010000e-07 V_low
+ 8.982000000e-07 V_low
+ 8.982010000e-07 V_low
+ 8.983000000e-07 V_low
+ 8.983010000e-07 V_low
+ 8.984000000e-07 V_low
+ 8.984010000e-07 V_low
+ 8.985000000e-07 V_low
+ 8.985010000e-07 V_low
+ 8.986000000e-07 V_low
+ 8.986010000e-07 V_low
+ 8.987000000e-07 V_low
+ 8.987010000e-07 V_low
+ 8.988000000e-07 V_low
+ 8.988010000e-07 V_low
+ 8.989000000e-07 V_low
+ 8.989010000e-07 V_low
+ 8.990000000e-07 V_low
+ 8.990010000e-07 V_low
+ 8.991000000e-07 V_low
+ 8.991010000e-07 V_low
+ 8.992000000e-07 V_low
+ 8.992010000e-07 V_low
+ 8.993000000e-07 V_low
+ 8.993010000e-07 V_low
+ 8.994000000e-07 V_low
+ 8.994010000e-07 V_low
+ 8.995000000e-07 V_low
+ 8.995010000e-07 V_low
+ 8.996000000e-07 V_low
+ 8.996010000e-07 V_low
+ 8.997000000e-07 V_low
+ 8.997010000e-07 V_low
+ 8.998000000e-07 V_low
+ 8.998010000e-07 V_low
+ 8.999000000e-07 V_low
+ 8.999010000e-07 V_low
+ 9.000000000e-07 V_low
+ 9.000010000e-07 V_low
+ 9.001000000e-07 V_low
+ 9.001010000e-07 V_low
+ 9.002000000e-07 V_low
+ 9.002010000e-07 V_low
+ 9.003000000e-07 V_low
+ 9.003010000e-07 V_low
+ 9.004000000e-07 V_low
+ 9.004010000e-07 V_low
+ 9.005000000e-07 V_low
+ 9.005010000e-07 V_low
+ 9.006000000e-07 V_low
+ 9.006010000e-07 V_low
+ 9.007000000e-07 V_low
+ 9.007010000e-07 V_low
+ 9.008000000e-07 V_low
+ 9.008010000e-07 V_low
+ 9.009000000e-07 V_low
+ 9.009010000e-07 V_low
+ 9.010000000e-07 V_low
+ 9.010010000e-07 V_low
+ 9.011000000e-07 V_low
+ 9.011010000e-07 V_low
+ 9.012000000e-07 V_low
+ 9.012010000e-07 V_low
+ 9.013000000e-07 V_low
+ 9.013010000e-07 V_low
+ 9.014000000e-07 V_low
+ 9.014010000e-07 V_low
+ 9.015000000e-07 V_low
+ 9.015010000e-07 V_low
+ 9.016000000e-07 V_low
+ 9.016010000e-07 V_low
+ 9.017000000e-07 V_low
+ 9.017010000e-07 V_low
+ 9.018000000e-07 V_low
+ 9.018010000e-07 V_low
+ 9.019000000e-07 V_low
+ 9.019010000e-07 V_low
+ 9.020000000e-07 V_low
+ 9.020010000e-07 V_low
+ 9.021000000e-07 V_low
+ 9.021010000e-07 V_low
+ 9.022000000e-07 V_low
+ 9.022010000e-07 V_low
+ 9.023000000e-07 V_low
+ 9.023010000e-07 V_low
+ 9.024000000e-07 V_low
+ 9.024010000e-07 V_low
+ 9.025000000e-07 V_low
+ 9.025010000e-07 V_low
+ 9.026000000e-07 V_low
+ 9.026010000e-07 V_low
+ 9.027000000e-07 V_low
+ 9.027010000e-07 V_low
+ 9.028000000e-07 V_low
+ 9.028010000e-07 V_low
+ 9.029000000e-07 V_low
+ 9.029010000e-07 V_hig
+ 9.030000000e-07 V_hig
+ 9.030010000e-07 V_hig
+ 9.031000000e-07 V_hig
+ 9.031010000e-07 V_hig
+ 9.032000000e-07 V_hig
+ 9.032010000e-07 V_hig
+ 9.033000000e-07 V_hig
+ 9.033010000e-07 V_hig
+ 9.034000000e-07 V_hig
+ 9.034010000e-07 V_hig
+ 9.035000000e-07 V_hig
+ 9.035010000e-07 V_hig
+ 9.036000000e-07 V_hig
+ 9.036010000e-07 V_hig
+ 9.037000000e-07 V_hig
+ 9.037010000e-07 V_hig
+ 9.038000000e-07 V_hig
+ 9.038010000e-07 V_hig
+ 9.039000000e-07 V_hig
+ 9.039010000e-07 V_hig
+ 9.040000000e-07 V_hig
+ 9.040010000e-07 V_hig
+ 9.041000000e-07 V_hig
+ 9.041010000e-07 V_hig
+ 9.042000000e-07 V_hig
+ 9.042010000e-07 V_hig
+ 9.043000000e-07 V_hig
+ 9.043010000e-07 V_hig
+ 9.044000000e-07 V_hig
+ 9.044010000e-07 V_hig
+ 9.045000000e-07 V_hig
+ 9.045010000e-07 V_hig
+ 9.046000000e-07 V_hig
+ 9.046010000e-07 V_hig
+ 9.047000000e-07 V_hig
+ 9.047010000e-07 V_hig
+ 9.048000000e-07 V_hig
+ 9.048010000e-07 V_hig
+ 9.049000000e-07 V_hig
+ 9.049010000e-07 V_hig
+ 9.050000000e-07 V_hig
+ 9.050010000e-07 V_hig
+ 9.051000000e-07 V_hig
+ 9.051010000e-07 V_hig
+ 9.052000000e-07 V_hig
+ 9.052010000e-07 V_hig
+ 9.053000000e-07 V_hig
+ 9.053010000e-07 V_hig
+ 9.054000000e-07 V_hig
+ 9.054010000e-07 V_hig
+ 9.055000000e-07 V_hig
+ 9.055010000e-07 V_hig
+ 9.056000000e-07 V_hig
+ 9.056010000e-07 V_hig
+ 9.057000000e-07 V_hig
+ 9.057010000e-07 V_hig
+ 9.058000000e-07 V_hig
+ 9.058010000e-07 V_hig
+ 9.059000000e-07 V_hig
+ 9.059010000e-07 V_low
+ 9.060000000e-07 V_low
+ 9.060010000e-07 V_low
+ 9.061000000e-07 V_low
+ 9.061010000e-07 V_low
+ 9.062000000e-07 V_low
+ 9.062010000e-07 V_low
+ 9.063000000e-07 V_low
+ 9.063010000e-07 V_low
+ 9.064000000e-07 V_low
+ 9.064010000e-07 V_low
+ 9.065000000e-07 V_low
+ 9.065010000e-07 V_low
+ 9.066000000e-07 V_low
+ 9.066010000e-07 V_low
+ 9.067000000e-07 V_low
+ 9.067010000e-07 V_low
+ 9.068000000e-07 V_low
+ 9.068010000e-07 V_low
+ 9.069000000e-07 V_low
+ 9.069010000e-07 V_hig
+ 9.070000000e-07 V_hig
+ 9.070010000e-07 V_hig
+ 9.071000000e-07 V_hig
+ 9.071010000e-07 V_hig
+ 9.072000000e-07 V_hig
+ 9.072010000e-07 V_hig
+ 9.073000000e-07 V_hig
+ 9.073010000e-07 V_hig
+ 9.074000000e-07 V_hig
+ 9.074010000e-07 V_hig
+ 9.075000000e-07 V_hig
+ 9.075010000e-07 V_hig
+ 9.076000000e-07 V_hig
+ 9.076010000e-07 V_hig
+ 9.077000000e-07 V_hig
+ 9.077010000e-07 V_hig
+ 9.078000000e-07 V_hig
+ 9.078010000e-07 V_hig
+ 9.079000000e-07 V_hig
+ 9.079010000e-07 V_hig
+ 9.080000000e-07 V_hig
+ 9.080010000e-07 V_hig
+ 9.081000000e-07 V_hig
+ 9.081010000e-07 V_hig
+ 9.082000000e-07 V_hig
+ 9.082010000e-07 V_hig
+ 9.083000000e-07 V_hig
+ 9.083010000e-07 V_hig
+ 9.084000000e-07 V_hig
+ 9.084010000e-07 V_hig
+ 9.085000000e-07 V_hig
+ 9.085010000e-07 V_hig
+ 9.086000000e-07 V_hig
+ 9.086010000e-07 V_hig
+ 9.087000000e-07 V_hig
+ 9.087010000e-07 V_hig
+ 9.088000000e-07 V_hig
+ 9.088010000e-07 V_hig
+ 9.089000000e-07 V_hig
+ 9.089010000e-07 V_low
+ 9.090000000e-07 V_low
+ 9.090010000e-07 V_low
+ 9.091000000e-07 V_low
+ 9.091010000e-07 V_low
+ 9.092000000e-07 V_low
+ 9.092010000e-07 V_low
+ 9.093000000e-07 V_low
+ 9.093010000e-07 V_low
+ 9.094000000e-07 V_low
+ 9.094010000e-07 V_low
+ 9.095000000e-07 V_low
+ 9.095010000e-07 V_low
+ 9.096000000e-07 V_low
+ 9.096010000e-07 V_low
+ 9.097000000e-07 V_low
+ 9.097010000e-07 V_low
+ 9.098000000e-07 V_low
+ 9.098010000e-07 V_low
+ 9.099000000e-07 V_low
+ 9.099010000e-07 V_low
+ 9.100000000e-07 V_low
+ 9.100010000e-07 V_low
+ 9.101000000e-07 V_low
+ 9.101010000e-07 V_low
+ 9.102000000e-07 V_low
+ 9.102010000e-07 V_low
+ 9.103000000e-07 V_low
+ 9.103010000e-07 V_low
+ 9.104000000e-07 V_low
+ 9.104010000e-07 V_low
+ 9.105000000e-07 V_low
+ 9.105010000e-07 V_low
+ 9.106000000e-07 V_low
+ 9.106010000e-07 V_low
+ 9.107000000e-07 V_low
+ 9.107010000e-07 V_low
+ 9.108000000e-07 V_low
+ 9.108010000e-07 V_low
+ 9.109000000e-07 V_low
+ 9.109010000e-07 V_low
+ 9.110000000e-07 V_low
+ 9.110010000e-07 V_low
+ 9.111000000e-07 V_low
+ 9.111010000e-07 V_low
+ 9.112000000e-07 V_low
+ 9.112010000e-07 V_low
+ 9.113000000e-07 V_low
+ 9.113010000e-07 V_low
+ 9.114000000e-07 V_low
+ 9.114010000e-07 V_low
+ 9.115000000e-07 V_low
+ 9.115010000e-07 V_low
+ 9.116000000e-07 V_low
+ 9.116010000e-07 V_low
+ 9.117000000e-07 V_low
+ 9.117010000e-07 V_low
+ 9.118000000e-07 V_low
+ 9.118010000e-07 V_low
+ 9.119000000e-07 V_low
+ 9.119010000e-07 V_low
+ 9.120000000e-07 V_low
+ 9.120010000e-07 V_low
+ 9.121000000e-07 V_low
+ 9.121010000e-07 V_low
+ 9.122000000e-07 V_low
+ 9.122010000e-07 V_low
+ 9.123000000e-07 V_low
+ 9.123010000e-07 V_low
+ 9.124000000e-07 V_low
+ 9.124010000e-07 V_low
+ 9.125000000e-07 V_low
+ 9.125010000e-07 V_low
+ 9.126000000e-07 V_low
+ 9.126010000e-07 V_low
+ 9.127000000e-07 V_low
+ 9.127010000e-07 V_low
+ 9.128000000e-07 V_low
+ 9.128010000e-07 V_low
+ 9.129000000e-07 V_low
+ 9.129010000e-07 V_hig
+ 9.130000000e-07 V_hig
+ 9.130010000e-07 V_hig
+ 9.131000000e-07 V_hig
+ 9.131010000e-07 V_hig
+ 9.132000000e-07 V_hig
+ 9.132010000e-07 V_hig
+ 9.133000000e-07 V_hig
+ 9.133010000e-07 V_hig
+ 9.134000000e-07 V_hig
+ 9.134010000e-07 V_hig
+ 9.135000000e-07 V_hig
+ 9.135010000e-07 V_hig
+ 9.136000000e-07 V_hig
+ 9.136010000e-07 V_hig
+ 9.137000000e-07 V_hig
+ 9.137010000e-07 V_hig
+ 9.138000000e-07 V_hig
+ 9.138010000e-07 V_hig
+ 9.139000000e-07 V_hig
+ 9.139010000e-07 V_hig
+ 9.140000000e-07 V_hig
+ 9.140010000e-07 V_hig
+ 9.141000000e-07 V_hig
+ 9.141010000e-07 V_hig
+ 9.142000000e-07 V_hig
+ 9.142010000e-07 V_hig
+ 9.143000000e-07 V_hig
+ 9.143010000e-07 V_hig
+ 9.144000000e-07 V_hig
+ 9.144010000e-07 V_hig
+ 9.145000000e-07 V_hig
+ 9.145010000e-07 V_hig
+ 9.146000000e-07 V_hig
+ 9.146010000e-07 V_hig
+ 9.147000000e-07 V_hig
+ 9.147010000e-07 V_hig
+ 9.148000000e-07 V_hig
+ 9.148010000e-07 V_hig
+ 9.149000000e-07 V_hig
+ 9.149010000e-07 V_low
+ 9.150000000e-07 V_low
+ 9.150010000e-07 V_low
+ 9.151000000e-07 V_low
+ 9.151010000e-07 V_low
+ 9.152000000e-07 V_low
+ 9.152010000e-07 V_low
+ 9.153000000e-07 V_low
+ 9.153010000e-07 V_low
+ 9.154000000e-07 V_low
+ 9.154010000e-07 V_low
+ 9.155000000e-07 V_low
+ 9.155010000e-07 V_low
+ 9.156000000e-07 V_low
+ 9.156010000e-07 V_low
+ 9.157000000e-07 V_low
+ 9.157010000e-07 V_low
+ 9.158000000e-07 V_low
+ 9.158010000e-07 V_low
+ 9.159000000e-07 V_low
+ 9.159010000e-07 V_hig
+ 9.160000000e-07 V_hig
+ 9.160010000e-07 V_hig
+ 9.161000000e-07 V_hig
+ 9.161010000e-07 V_hig
+ 9.162000000e-07 V_hig
+ 9.162010000e-07 V_hig
+ 9.163000000e-07 V_hig
+ 9.163010000e-07 V_hig
+ 9.164000000e-07 V_hig
+ 9.164010000e-07 V_hig
+ 9.165000000e-07 V_hig
+ 9.165010000e-07 V_hig
+ 9.166000000e-07 V_hig
+ 9.166010000e-07 V_hig
+ 9.167000000e-07 V_hig
+ 9.167010000e-07 V_hig
+ 9.168000000e-07 V_hig
+ 9.168010000e-07 V_hig
+ 9.169000000e-07 V_hig
+ 9.169010000e-07 V_low
+ 9.170000000e-07 V_low
+ 9.170010000e-07 V_low
+ 9.171000000e-07 V_low
+ 9.171010000e-07 V_low
+ 9.172000000e-07 V_low
+ 9.172010000e-07 V_low
+ 9.173000000e-07 V_low
+ 9.173010000e-07 V_low
+ 9.174000000e-07 V_low
+ 9.174010000e-07 V_low
+ 9.175000000e-07 V_low
+ 9.175010000e-07 V_low
+ 9.176000000e-07 V_low
+ 9.176010000e-07 V_low
+ 9.177000000e-07 V_low
+ 9.177010000e-07 V_low
+ 9.178000000e-07 V_low
+ 9.178010000e-07 V_low
+ 9.179000000e-07 V_low
+ 9.179010000e-07 V_low
+ 9.180000000e-07 V_low
+ 9.180010000e-07 V_low
+ 9.181000000e-07 V_low
+ 9.181010000e-07 V_low
+ 9.182000000e-07 V_low
+ 9.182010000e-07 V_low
+ 9.183000000e-07 V_low
+ 9.183010000e-07 V_low
+ 9.184000000e-07 V_low
+ 9.184010000e-07 V_low
+ 9.185000000e-07 V_low
+ 9.185010000e-07 V_low
+ 9.186000000e-07 V_low
+ 9.186010000e-07 V_low
+ 9.187000000e-07 V_low
+ 9.187010000e-07 V_low
+ 9.188000000e-07 V_low
+ 9.188010000e-07 V_low
+ 9.189000000e-07 V_low
+ 9.189010000e-07 V_low
+ 9.190000000e-07 V_low
+ 9.190010000e-07 V_low
+ 9.191000000e-07 V_low
+ 9.191010000e-07 V_low
+ 9.192000000e-07 V_low
+ 9.192010000e-07 V_low
+ 9.193000000e-07 V_low
+ 9.193010000e-07 V_low
+ 9.194000000e-07 V_low
+ 9.194010000e-07 V_low
+ 9.195000000e-07 V_low
+ 9.195010000e-07 V_low
+ 9.196000000e-07 V_low
+ 9.196010000e-07 V_low
+ 9.197000000e-07 V_low
+ 9.197010000e-07 V_low
+ 9.198000000e-07 V_low
+ 9.198010000e-07 V_low
+ 9.199000000e-07 V_low
+ 9.199010000e-07 V_low
+ 9.200000000e-07 V_low
+ 9.200010000e-07 V_low
+ 9.201000000e-07 V_low
+ 9.201010000e-07 V_low
+ 9.202000000e-07 V_low
+ 9.202010000e-07 V_low
+ 9.203000000e-07 V_low
+ 9.203010000e-07 V_low
+ 9.204000000e-07 V_low
+ 9.204010000e-07 V_low
+ 9.205000000e-07 V_low
+ 9.205010000e-07 V_low
+ 9.206000000e-07 V_low
+ 9.206010000e-07 V_low
+ 9.207000000e-07 V_low
+ 9.207010000e-07 V_low
+ 9.208000000e-07 V_low
+ 9.208010000e-07 V_low
+ 9.209000000e-07 V_low
+ 9.209010000e-07 V_hig
+ 9.210000000e-07 V_hig
+ 9.210010000e-07 V_hig
+ 9.211000000e-07 V_hig
+ 9.211010000e-07 V_hig
+ 9.212000000e-07 V_hig
+ 9.212010000e-07 V_hig
+ 9.213000000e-07 V_hig
+ 9.213010000e-07 V_hig
+ 9.214000000e-07 V_hig
+ 9.214010000e-07 V_hig
+ 9.215000000e-07 V_hig
+ 9.215010000e-07 V_hig
+ 9.216000000e-07 V_hig
+ 9.216010000e-07 V_hig
+ 9.217000000e-07 V_hig
+ 9.217010000e-07 V_hig
+ 9.218000000e-07 V_hig
+ 9.218010000e-07 V_hig
+ 9.219000000e-07 V_hig
+ 9.219010000e-07 V_hig
+ 9.220000000e-07 V_hig
+ 9.220010000e-07 V_hig
+ 9.221000000e-07 V_hig
+ 9.221010000e-07 V_hig
+ 9.222000000e-07 V_hig
+ 9.222010000e-07 V_hig
+ 9.223000000e-07 V_hig
+ 9.223010000e-07 V_hig
+ 9.224000000e-07 V_hig
+ 9.224010000e-07 V_hig
+ 9.225000000e-07 V_hig
+ 9.225010000e-07 V_hig
+ 9.226000000e-07 V_hig
+ 9.226010000e-07 V_hig
+ 9.227000000e-07 V_hig
+ 9.227010000e-07 V_hig
+ 9.228000000e-07 V_hig
+ 9.228010000e-07 V_hig
+ 9.229000000e-07 V_hig
+ 9.229010000e-07 V_low
+ 9.230000000e-07 V_low
+ 9.230010000e-07 V_low
+ 9.231000000e-07 V_low
+ 9.231010000e-07 V_low
+ 9.232000000e-07 V_low
+ 9.232010000e-07 V_low
+ 9.233000000e-07 V_low
+ 9.233010000e-07 V_low
+ 9.234000000e-07 V_low
+ 9.234010000e-07 V_low
+ 9.235000000e-07 V_low
+ 9.235010000e-07 V_low
+ 9.236000000e-07 V_low
+ 9.236010000e-07 V_low
+ 9.237000000e-07 V_low
+ 9.237010000e-07 V_low
+ 9.238000000e-07 V_low
+ 9.238010000e-07 V_low
+ 9.239000000e-07 V_low
+ 9.239010000e-07 V_low
+ 9.240000000e-07 V_low
+ 9.240010000e-07 V_low
+ 9.241000000e-07 V_low
+ 9.241010000e-07 V_low
+ 9.242000000e-07 V_low
+ 9.242010000e-07 V_low
+ 9.243000000e-07 V_low
+ 9.243010000e-07 V_low
+ 9.244000000e-07 V_low
+ 9.244010000e-07 V_low
+ 9.245000000e-07 V_low
+ 9.245010000e-07 V_low
+ 9.246000000e-07 V_low
+ 9.246010000e-07 V_low
+ 9.247000000e-07 V_low
+ 9.247010000e-07 V_low
+ 9.248000000e-07 V_low
+ 9.248010000e-07 V_low
+ 9.249000000e-07 V_low
+ 9.249010000e-07 V_low
+ 9.250000000e-07 V_low
+ 9.250010000e-07 V_low
+ 9.251000000e-07 V_low
+ 9.251010000e-07 V_low
+ 9.252000000e-07 V_low
+ 9.252010000e-07 V_low
+ 9.253000000e-07 V_low
+ 9.253010000e-07 V_low
+ 9.254000000e-07 V_low
+ 9.254010000e-07 V_low
+ 9.255000000e-07 V_low
+ 9.255010000e-07 V_low
+ 9.256000000e-07 V_low
+ 9.256010000e-07 V_low
+ 9.257000000e-07 V_low
+ 9.257010000e-07 V_low
+ 9.258000000e-07 V_low
+ 9.258010000e-07 V_low
+ 9.259000000e-07 V_low
+ 9.259010000e-07 V_low
+ 9.260000000e-07 V_low
+ 9.260010000e-07 V_low
+ 9.261000000e-07 V_low
+ 9.261010000e-07 V_low
+ 9.262000000e-07 V_low
+ 9.262010000e-07 V_low
+ 9.263000000e-07 V_low
+ 9.263010000e-07 V_low
+ 9.264000000e-07 V_low
+ 9.264010000e-07 V_low
+ 9.265000000e-07 V_low
+ 9.265010000e-07 V_low
+ 9.266000000e-07 V_low
+ 9.266010000e-07 V_low
+ 9.267000000e-07 V_low
+ 9.267010000e-07 V_low
+ 9.268000000e-07 V_low
+ 9.268010000e-07 V_low
+ 9.269000000e-07 V_low
+ 9.269010000e-07 V_hig
+ 9.270000000e-07 V_hig
+ 9.270010000e-07 V_hig
+ 9.271000000e-07 V_hig
+ 9.271010000e-07 V_hig
+ 9.272000000e-07 V_hig
+ 9.272010000e-07 V_hig
+ 9.273000000e-07 V_hig
+ 9.273010000e-07 V_hig
+ 9.274000000e-07 V_hig
+ 9.274010000e-07 V_hig
+ 9.275000000e-07 V_hig
+ 9.275010000e-07 V_hig
+ 9.276000000e-07 V_hig
+ 9.276010000e-07 V_hig
+ 9.277000000e-07 V_hig
+ 9.277010000e-07 V_hig
+ 9.278000000e-07 V_hig
+ 9.278010000e-07 V_hig
+ 9.279000000e-07 V_hig
+ 9.279010000e-07 V_low
+ 9.280000000e-07 V_low
+ 9.280010000e-07 V_low
+ 9.281000000e-07 V_low
+ 9.281010000e-07 V_low
+ 9.282000000e-07 V_low
+ 9.282010000e-07 V_low
+ 9.283000000e-07 V_low
+ 9.283010000e-07 V_low
+ 9.284000000e-07 V_low
+ 9.284010000e-07 V_low
+ 9.285000000e-07 V_low
+ 9.285010000e-07 V_low
+ 9.286000000e-07 V_low
+ 9.286010000e-07 V_low
+ 9.287000000e-07 V_low
+ 9.287010000e-07 V_low
+ 9.288000000e-07 V_low
+ 9.288010000e-07 V_low
+ 9.289000000e-07 V_low
+ 9.289010000e-07 V_low
+ 9.290000000e-07 V_low
+ 9.290010000e-07 V_low
+ 9.291000000e-07 V_low
+ 9.291010000e-07 V_low
+ 9.292000000e-07 V_low
+ 9.292010000e-07 V_low
+ 9.293000000e-07 V_low
+ 9.293010000e-07 V_low
+ 9.294000000e-07 V_low
+ 9.294010000e-07 V_low
+ 9.295000000e-07 V_low
+ 9.295010000e-07 V_low
+ 9.296000000e-07 V_low
+ 9.296010000e-07 V_low
+ 9.297000000e-07 V_low
+ 9.297010000e-07 V_low
+ 9.298000000e-07 V_low
+ 9.298010000e-07 V_low
+ 9.299000000e-07 V_low
+ 9.299010000e-07 V_hig
+ 9.300000000e-07 V_hig
+ 9.300010000e-07 V_hig
+ 9.301000000e-07 V_hig
+ 9.301010000e-07 V_hig
+ 9.302000000e-07 V_hig
+ 9.302010000e-07 V_hig
+ 9.303000000e-07 V_hig
+ 9.303010000e-07 V_hig
+ 9.304000000e-07 V_hig
+ 9.304010000e-07 V_hig
+ 9.305000000e-07 V_hig
+ 9.305010000e-07 V_hig
+ 9.306000000e-07 V_hig
+ 9.306010000e-07 V_hig
+ 9.307000000e-07 V_hig
+ 9.307010000e-07 V_hig
+ 9.308000000e-07 V_hig
+ 9.308010000e-07 V_hig
+ 9.309000000e-07 V_hig
+ 9.309010000e-07 V_hig
+ 9.310000000e-07 V_hig
+ 9.310010000e-07 V_hig
+ 9.311000000e-07 V_hig
+ 9.311010000e-07 V_hig
+ 9.312000000e-07 V_hig
+ 9.312010000e-07 V_hig
+ 9.313000000e-07 V_hig
+ 9.313010000e-07 V_hig
+ 9.314000000e-07 V_hig
+ 9.314010000e-07 V_hig
+ 9.315000000e-07 V_hig
+ 9.315010000e-07 V_hig
+ 9.316000000e-07 V_hig
+ 9.316010000e-07 V_hig
+ 9.317000000e-07 V_hig
+ 9.317010000e-07 V_hig
+ 9.318000000e-07 V_hig
+ 9.318010000e-07 V_hig
+ 9.319000000e-07 V_hig
+ 9.319010000e-07 V_hig
+ 9.320000000e-07 V_hig
+ 9.320010000e-07 V_hig
+ 9.321000000e-07 V_hig
+ 9.321010000e-07 V_hig
+ 9.322000000e-07 V_hig
+ 9.322010000e-07 V_hig
+ 9.323000000e-07 V_hig
+ 9.323010000e-07 V_hig
+ 9.324000000e-07 V_hig
+ 9.324010000e-07 V_hig
+ 9.325000000e-07 V_hig
+ 9.325010000e-07 V_hig
+ 9.326000000e-07 V_hig
+ 9.326010000e-07 V_hig
+ 9.327000000e-07 V_hig
+ 9.327010000e-07 V_hig
+ 9.328000000e-07 V_hig
+ 9.328010000e-07 V_hig
+ 9.329000000e-07 V_hig
+ 9.329010000e-07 V_hig
+ 9.330000000e-07 V_hig
+ 9.330010000e-07 V_hig
+ 9.331000000e-07 V_hig
+ 9.331010000e-07 V_hig
+ 9.332000000e-07 V_hig
+ 9.332010000e-07 V_hig
+ 9.333000000e-07 V_hig
+ 9.333010000e-07 V_hig
+ 9.334000000e-07 V_hig
+ 9.334010000e-07 V_hig
+ 9.335000000e-07 V_hig
+ 9.335010000e-07 V_hig
+ 9.336000000e-07 V_hig
+ 9.336010000e-07 V_hig
+ 9.337000000e-07 V_hig
+ 9.337010000e-07 V_hig
+ 9.338000000e-07 V_hig
+ 9.338010000e-07 V_hig
+ 9.339000000e-07 V_hig
+ 9.339010000e-07 V_hig
+ 9.340000000e-07 V_hig
+ 9.340010000e-07 V_hig
+ 9.341000000e-07 V_hig
+ 9.341010000e-07 V_hig
+ 9.342000000e-07 V_hig
+ 9.342010000e-07 V_hig
+ 9.343000000e-07 V_hig
+ 9.343010000e-07 V_hig
+ 9.344000000e-07 V_hig
+ 9.344010000e-07 V_hig
+ 9.345000000e-07 V_hig
+ 9.345010000e-07 V_hig
+ 9.346000000e-07 V_hig
+ 9.346010000e-07 V_hig
+ 9.347000000e-07 V_hig
+ 9.347010000e-07 V_hig
+ 9.348000000e-07 V_hig
+ 9.348010000e-07 V_hig
+ 9.349000000e-07 V_hig
+ 9.349010000e-07 V_hig
+ 9.350000000e-07 V_hig
+ 9.350010000e-07 V_hig
+ 9.351000000e-07 V_hig
+ 9.351010000e-07 V_hig
+ 9.352000000e-07 V_hig
+ 9.352010000e-07 V_hig
+ 9.353000000e-07 V_hig
+ 9.353010000e-07 V_hig
+ 9.354000000e-07 V_hig
+ 9.354010000e-07 V_hig
+ 9.355000000e-07 V_hig
+ 9.355010000e-07 V_hig
+ 9.356000000e-07 V_hig
+ 9.356010000e-07 V_hig
+ 9.357000000e-07 V_hig
+ 9.357010000e-07 V_hig
+ 9.358000000e-07 V_hig
+ 9.358010000e-07 V_hig
+ 9.359000000e-07 V_hig
+ 9.359010000e-07 V_hig
+ 9.360000000e-07 V_hig
+ 9.360010000e-07 V_hig
+ 9.361000000e-07 V_hig
+ 9.361010000e-07 V_hig
+ 9.362000000e-07 V_hig
+ 9.362010000e-07 V_hig
+ 9.363000000e-07 V_hig
+ 9.363010000e-07 V_hig
+ 9.364000000e-07 V_hig
+ 9.364010000e-07 V_hig
+ 9.365000000e-07 V_hig
+ 9.365010000e-07 V_hig
+ 9.366000000e-07 V_hig
+ 9.366010000e-07 V_hig
+ 9.367000000e-07 V_hig
+ 9.367010000e-07 V_hig
+ 9.368000000e-07 V_hig
+ 9.368010000e-07 V_hig
+ 9.369000000e-07 V_hig
+ 9.369010000e-07 V_low
+ 9.370000000e-07 V_low
+ 9.370010000e-07 V_low
+ 9.371000000e-07 V_low
+ 9.371010000e-07 V_low
+ 9.372000000e-07 V_low
+ 9.372010000e-07 V_low
+ 9.373000000e-07 V_low
+ 9.373010000e-07 V_low
+ 9.374000000e-07 V_low
+ 9.374010000e-07 V_low
+ 9.375000000e-07 V_low
+ 9.375010000e-07 V_low
+ 9.376000000e-07 V_low
+ 9.376010000e-07 V_low
+ 9.377000000e-07 V_low
+ 9.377010000e-07 V_low
+ 9.378000000e-07 V_low
+ 9.378010000e-07 V_low
+ 9.379000000e-07 V_low
+ 9.379010000e-07 V_hig
+ 9.380000000e-07 V_hig
+ 9.380010000e-07 V_hig
+ 9.381000000e-07 V_hig
+ 9.381010000e-07 V_hig
+ 9.382000000e-07 V_hig
+ 9.382010000e-07 V_hig
+ 9.383000000e-07 V_hig
+ 9.383010000e-07 V_hig
+ 9.384000000e-07 V_hig
+ 9.384010000e-07 V_hig
+ 9.385000000e-07 V_hig
+ 9.385010000e-07 V_hig
+ 9.386000000e-07 V_hig
+ 9.386010000e-07 V_hig
+ 9.387000000e-07 V_hig
+ 9.387010000e-07 V_hig
+ 9.388000000e-07 V_hig
+ 9.388010000e-07 V_hig
+ 9.389000000e-07 V_hig
+ 9.389010000e-07 V_low
+ 9.390000000e-07 V_low
+ 9.390010000e-07 V_low
+ 9.391000000e-07 V_low
+ 9.391010000e-07 V_low
+ 9.392000000e-07 V_low
+ 9.392010000e-07 V_low
+ 9.393000000e-07 V_low
+ 9.393010000e-07 V_low
+ 9.394000000e-07 V_low
+ 9.394010000e-07 V_low
+ 9.395000000e-07 V_low
+ 9.395010000e-07 V_low
+ 9.396000000e-07 V_low
+ 9.396010000e-07 V_low
+ 9.397000000e-07 V_low
+ 9.397010000e-07 V_low
+ 9.398000000e-07 V_low
+ 9.398010000e-07 V_low
+ 9.399000000e-07 V_low
+ 9.399010000e-07 V_hig
+ 9.400000000e-07 V_hig
+ 9.400010000e-07 V_hig
+ 9.401000000e-07 V_hig
+ 9.401010000e-07 V_hig
+ 9.402000000e-07 V_hig
+ 9.402010000e-07 V_hig
+ 9.403000000e-07 V_hig
+ 9.403010000e-07 V_hig
+ 9.404000000e-07 V_hig
+ 9.404010000e-07 V_hig
+ 9.405000000e-07 V_hig
+ 9.405010000e-07 V_hig
+ 9.406000000e-07 V_hig
+ 9.406010000e-07 V_hig
+ 9.407000000e-07 V_hig
+ 9.407010000e-07 V_hig
+ 9.408000000e-07 V_hig
+ 9.408010000e-07 V_hig
+ 9.409000000e-07 V_hig
+ 9.409010000e-07 V_low
+ 9.410000000e-07 V_low
+ 9.410010000e-07 V_low
+ 9.411000000e-07 V_low
+ 9.411010000e-07 V_low
+ 9.412000000e-07 V_low
+ 9.412010000e-07 V_low
+ 9.413000000e-07 V_low
+ 9.413010000e-07 V_low
+ 9.414000000e-07 V_low
+ 9.414010000e-07 V_low
+ 9.415000000e-07 V_low
+ 9.415010000e-07 V_low
+ 9.416000000e-07 V_low
+ 9.416010000e-07 V_low
+ 9.417000000e-07 V_low
+ 9.417010000e-07 V_low
+ 9.418000000e-07 V_low
+ 9.418010000e-07 V_low
+ 9.419000000e-07 V_low
+ 9.419010000e-07 V_low
+ 9.420000000e-07 V_low
+ 9.420010000e-07 V_low
+ 9.421000000e-07 V_low
+ 9.421010000e-07 V_low
+ 9.422000000e-07 V_low
+ 9.422010000e-07 V_low
+ 9.423000000e-07 V_low
+ 9.423010000e-07 V_low
+ 9.424000000e-07 V_low
+ 9.424010000e-07 V_low
+ 9.425000000e-07 V_low
+ 9.425010000e-07 V_low
+ 9.426000000e-07 V_low
+ 9.426010000e-07 V_low
+ 9.427000000e-07 V_low
+ 9.427010000e-07 V_low
+ 9.428000000e-07 V_low
+ 9.428010000e-07 V_low
+ 9.429000000e-07 V_low
+ 9.429010000e-07 V_low
+ 9.430000000e-07 V_low
+ 9.430010000e-07 V_low
+ 9.431000000e-07 V_low
+ 9.431010000e-07 V_low
+ 9.432000000e-07 V_low
+ 9.432010000e-07 V_low
+ 9.433000000e-07 V_low
+ 9.433010000e-07 V_low
+ 9.434000000e-07 V_low
+ 9.434010000e-07 V_low
+ 9.435000000e-07 V_low
+ 9.435010000e-07 V_low
+ 9.436000000e-07 V_low
+ 9.436010000e-07 V_low
+ 9.437000000e-07 V_low
+ 9.437010000e-07 V_low
+ 9.438000000e-07 V_low
+ 9.438010000e-07 V_low
+ 9.439000000e-07 V_low
+ 9.439010000e-07 V_low
+ 9.440000000e-07 V_low
+ 9.440010000e-07 V_low
+ 9.441000000e-07 V_low
+ 9.441010000e-07 V_low
+ 9.442000000e-07 V_low
+ 9.442010000e-07 V_low
+ 9.443000000e-07 V_low
+ 9.443010000e-07 V_low
+ 9.444000000e-07 V_low
+ 9.444010000e-07 V_low
+ 9.445000000e-07 V_low
+ 9.445010000e-07 V_low
+ 9.446000000e-07 V_low
+ 9.446010000e-07 V_low
+ 9.447000000e-07 V_low
+ 9.447010000e-07 V_low
+ 9.448000000e-07 V_low
+ 9.448010000e-07 V_low
+ 9.449000000e-07 V_low
+ 9.449010000e-07 V_low
+ 9.450000000e-07 V_low
+ 9.450010000e-07 V_low
+ 9.451000000e-07 V_low
+ 9.451010000e-07 V_low
+ 9.452000000e-07 V_low
+ 9.452010000e-07 V_low
+ 9.453000000e-07 V_low
+ 9.453010000e-07 V_low
+ 9.454000000e-07 V_low
+ 9.454010000e-07 V_low
+ 9.455000000e-07 V_low
+ 9.455010000e-07 V_low
+ 9.456000000e-07 V_low
+ 9.456010000e-07 V_low
+ 9.457000000e-07 V_low
+ 9.457010000e-07 V_low
+ 9.458000000e-07 V_low
+ 9.458010000e-07 V_low
+ 9.459000000e-07 V_low
+ 9.459010000e-07 V_low
+ 9.460000000e-07 V_low
+ 9.460010000e-07 V_low
+ 9.461000000e-07 V_low
+ 9.461010000e-07 V_low
+ 9.462000000e-07 V_low
+ 9.462010000e-07 V_low
+ 9.463000000e-07 V_low
+ 9.463010000e-07 V_low
+ 9.464000000e-07 V_low
+ 9.464010000e-07 V_low
+ 9.465000000e-07 V_low
+ 9.465010000e-07 V_low
+ 9.466000000e-07 V_low
+ 9.466010000e-07 V_low
+ 9.467000000e-07 V_low
+ 9.467010000e-07 V_low
+ 9.468000000e-07 V_low
+ 9.468010000e-07 V_low
+ 9.469000000e-07 V_low
+ 9.469010000e-07 V_hig
+ 9.470000000e-07 V_hig
+ 9.470010000e-07 V_hig
+ 9.471000000e-07 V_hig
+ 9.471010000e-07 V_hig
+ 9.472000000e-07 V_hig
+ 9.472010000e-07 V_hig
+ 9.473000000e-07 V_hig
+ 9.473010000e-07 V_hig
+ 9.474000000e-07 V_hig
+ 9.474010000e-07 V_hig
+ 9.475000000e-07 V_hig
+ 9.475010000e-07 V_hig
+ 9.476000000e-07 V_hig
+ 9.476010000e-07 V_hig
+ 9.477000000e-07 V_hig
+ 9.477010000e-07 V_hig
+ 9.478000000e-07 V_hig
+ 9.478010000e-07 V_hig
+ 9.479000000e-07 V_hig
+ 9.479010000e-07 V_hig
+ 9.480000000e-07 V_hig
+ 9.480010000e-07 V_hig
+ 9.481000000e-07 V_hig
+ 9.481010000e-07 V_hig
+ 9.482000000e-07 V_hig
+ 9.482010000e-07 V_hig
+ 9.483000000e-07 V_hig
+ 9.483010000e-07 V_hig
+ 9.484000000e-07 V_hig
+ 9.484010000e-07 V_hig
+ 9.485000000e-07 V_hig
+ 9.485010000e-07 V_hig
+ 9.486000000e-07 V_hig
+ 9.486010000e-07 V_hig
+ 9.487000000e-07 V_hig
+ 9.487010000e-07 V_hig
+ 9.488000000e-07 V_hig
+ 9.488010000e-07 V_hig
+ 9.489000000e-07 V_hig
+ 9.489010000e-07 V_hig
+ 9.490000000e-07 V_hig
+ 9.490010000e-07 V_hig
+ 9.491000000e-07 V_hig
+ 9.491010000e-07 V_hig
+ 9.492000000e-07 V_hig
+ 9.492010000e-07 V_hig
+ 9.493000000e-07 V_hig
+ 9.493010000e-07 V_hig
+ 9.494000000e-07 V_hig
+ 9.494010000e-07 V_hig
+ 9.495000000e-07 V_hig
+ 9.495010000e-07 V_hig
+ 9.496000000e-07 V_hig
+ 9.496010000e-07 V_hig
+ 9.497000000e-07 V_hig
+ 9.497010000e-07 V_hig
+ 9.498000000e-07 V_hig
+ 9.498010000e-07 V_hig
+ 9.499000000e-07 V_hig
+ 9.499010000e-07 V_low
+ 9.500000000e-07 V_low
+ 9.500010000e-07 V_low
+ 9.501000000e-07 V_low
+ 9.501010000e-07 V_low
+ 9.502000000e-07 V_low
+ 9.502010000e-07 V_low
+ 9.503000000e-07 V_low
+ 9.503010000e-07 V_low
+ 9.504000000e-07 V_low
+ 9.504010000e-07 V_low
+ 9.505000000e-07 V_low
+ 9.505010000e-07 V_low
+ 9.506000000e-07 V_low
+ 9.506010000e-07 V_low
+ 9.507000000e-07 V_low
+ 9.507010000e-07 V_low
+ 9.508000000e-07 V_low
+ 9.508010000e-07 V_low
+ 9.509000000e-07 V_low
+ 9.509010000e-07 V_hig
+ 9.510000000e-07 V_hig
+ 9.510010000e-07 V_hig
+ 9.511000000e-07 V_hig
+ 9.511010000e-07 V_hig
+ 9.512000000e-07 V_hig
+ 9.512010000e-07 V_hig
+ 9.513000000e-07 V_hig
+ 9.513010000e-07 V_hig
+ 9.514000000e-07 V_hig
+ 9.514010000e-07 V_hig
+ 9.515000000e-07 V_hig
+ 9.515010000e-07 V_hig
+ 9.516000000e-07 V_hig
+ 9.516010000e-07 V_hig
+ 9.517000000e-07 V_hig
+ 9.517010000e-07 V_hig
+ 9.518000000e-07 V_hig
+ 9.518010000e-07 V_hig
+ 9.519000000e-07 V_hig
+ 9.519010000e-07 V_low
+ 9.520000000e-07 V_low
+ 9.520010000e-07 V_low
+ 9.521000000e-07 V_low
+ 9.521010000e-07 V_low
+ 9.522000000e-07 V_low
+ 9.522010000e-07 V_low
+ 9.523000000e-07 V_low
+ 9.523010000e-07 V_low
+ 9.524000000e-07 V_low
+ 9.524010000e-07 V_low
+ 9.525000000e-07 V_low
+ 9.525010000e-07 V_low
+ 9.526000000e-07 V_low
+ 9.526010000e-07 V_low
+ 9.527000000e-07 V_low
+ 9.527010000e-07 V_low
+ 9.528000000e-07 V_low
+ 9.528010000e-07 V_low
+ 9.529000000e-07 V_low
+ 9.529010000e-07 V_low
+ 9.530000000e-07 V_low
+ 9.530010000e-07 V_low
+ 9.531000000e-07 V_low
+ 9.531010000e-07 V_low
+ 9.532000000e-07 V_low
+ 9.532010000e-07 V_low
+ 9.533000000e-07 V_low
+ 9.533010000e-07 V_low
+ 9.534000000e-07 V_low
+ 9.534010000e-07 V_low
+ 9.535000000e-07 V_low
+ 9.535010000e-07 V_low
+ 9.536000000e-07 V_low
+ 9.536010000e-07 V_low
+ 9.537000000e-07 V_low
+ 9.537010000e-07 V_low
+ 9.538000000e-07 V_low
+ 9.538010000e-07 V_low
+ 9.539000000e-07 V_low
+ 9.539010000e-07 V_low
+ 9.540000000e-07 V_low
+ 9.540010000e-07 V_low
+ 9.541000000e-07 V_low
+ 9.541010000e-07 V_low
+ 9.542000000e-07 V_low
+ 9.542010000e-07 V_low
+ 9.543000000e-07 V_low
+ 9.543010000e-07 V_low
+ 9.544000000e-07 V_low
+ 9.544010000e-07 V_low
+ 9.545000000e-07 V_low
+ 9.545010000e-07 V_low
+ 9.546000000e-07 V_low
+ 9.546010000e-07 V_low
+ 9.547000000e-07 V_low
+ 9.547010000e-07 V_low
+ 9.548000000e-07 V_low
+ 9.548010000e-07 V_low
+ 9.549000000e-07 V_low
+ 9.549010000e-07 V_low
+ 9.550000000e-07 V_low
+ 9.550010000e-07 V_low
+ 9.551000000e-07 V_low
+ 9.551010000e-07 V_low
+ 9.552000000e-07 V_low
+ 9.552010000e-07 V_low
+ 9.553000000e-07 V_low
+ 9.553010000e-07 V_low
+ 9.554000000e-07 V_low
+ 9.554010000e-07 V_low
+ 9.555000000e-07 V_low
+ 9.555010000e-07 V_low
+ 9.556000000e-07 V_low
+ 9.556010000e-07 V_low
+ 9.557000000e-07 V_low
+ 9.557010000e-07 V_low
+ 9.558000000e-07 V_low
+ 9.558010000e-07 V_low
+ 9.559000000e-07 V_low
+ 9.559010000e-07 V_hig
+ 9.560000000e-07 V_hig
+ 9.560010000e-07 V_hig
+ 9.561000000e-07 V_hig
+ 9.561010000e-07 V_hig
+ 9.562000000e-07 V_hig
+ 9.562010000e-07 V_hig
+ 9.563000000e-07 V_hig
+ 9.563010000e-07 V_hig
+ 9.564000000e-07 V_hig
+ 9.564010000e-07 V_hig
+ 9.565000000e-07 V_hig
+ 9.565010000e-07 V_hig
+ 9.566000000e-07 V_hig
+ 9.566010000e-07 V_hig
+ 9.567000000e-07 V_hig
+ 9.567010000e-07 V_hig
+ 9.568000000e-07 V_hig
+ 9.568010000e-07 V_hig
+ 9.569000000e-07 V_hig
+ 9.569010000e-07 V_low
+ 9.570000000e-07 V_low
+ 9.570010000e-07 V_low
+ 9.571000000e-07 V_low
+ 9.571010000e-07 V_low
+ 9.572000000e-07 V_low
+ 9.572010000e-07 V_low
+ 9.573000000e-07 V_low
+ 9.573010000e-07 V_low
+ 9.574000000e-07 V_low
+ 9.574010000e-07 V_low
+ 9.575000000e-07 V_low
+ 9.575010000e-07 V_low
+ 9.576000000e-07 V_low
+ 9.576010000e-07 V_low
+ 9.577000000e-07 V_low
+ 9.577010000e-07 V_low
+ 9.578000000e-07 V_low
+ 9.578010000e-07 V_low
+ 9.579000000e-07 V_low
+ 9.579010000e-07 V_low
+ 9.580000000e-07 V_low
+ 9.580010000e-07 V_low
+ 9.581000000e-07 V_low
+ 9.581010000e-07 V_low
+ 9.582000000e-07 V_low
+ 9.582010000e-07 V_low
+ 9.583000000e-07 V_low
+ 9.583010000e-07 V_low
+ 9.584000000e-07 V_low
+ 9.584010000e-07 V_low
+ 9.585000000e-07 V_low
+ 9.585010000e-07 V_low
+ 9.586000000e-07 V_low
+ 9.586010000e-07 V_low
+ 9.587000000e-07 V_low
+ 9.587010000e-07 V_low
+ 9.588000000e-07 V_low
+ 9.588010000e-07 V_low
+ 9.589000000e-07 V_low
+ 9.589010000e-07 V_hig
+ 9.590000000e-07 V_hig
+ 9.590010000e-07 V_hig
+ 9.591000000e-07 V_hig
+ 9.591010000e-07 V_hig
+ 9.592000000e-07 V_hig
+ 9.592010000e-07 V_hig
+ 9.593000000e-07 V_hig
+ 9.593010000e-07 V_hig
+ 9.594000000e-07 V_hig
+ 9.594010000e-07 V_hig
+ 9.595000000e-07 V_hig
+ 9.595010000e-07 V_hig
+ 9.596000000e-07 V_hig
+ 9.596010000e-07 V_hig
+ 9.597000000e-07 V_hig
+ 9.597010000e-07 V_hig
+ 9.598000000e-07 V_hig
+ 9.598010000e-07 V_hig
+ 9.599000000e-07 V_hig
+ 9.599010000e-07 V_hig
+ 9.600000000e-07 V_hig
+ 9.600010000e-07 V_hig
+ 9.601000000e-07 V_hig
+ 9.601010000e-07 V_hig
+ 9.602000000e-07 V_hig
+ 9.602010000e-07 V_hig
+ 9.603000000e-07 V_hig
+ 9.603010000e-07 V_hig
+ 9.604000000e-07 V_hig
+ 9.604010000e-07 V_hig
+ 9.605000000e-07 V_hig
+ 9.605010000e-07 V_hig
+ 9.606000000e-07 V_hig
+ 9.606010000e-07 V_hig
+ 9.607000000e-07 V_hig
+ 9.607010000e-07 V_hig
+ 9.608000000e-07 V_hig
+ 9.608010000e-07 V_hig
+ 9.609000000e-07 V_hig
+ 9.609010000e-07 V_low
+ 9.610000000e-07 V_low
+ 9.610010000e-07 V_low
+ 9.611000000e-07 V_low
+ 9.611010000e-07 V_low
+ 9.612000000e-07 V_low
+ 9.612010000e-07 V_low
+ 9.613000000e-07 V_low
+ 9.613010000e-07 V_low
+ 9.614000000e-07 V_low
+ 9.614010000e-07 V_low
+ 9.615000000e-07 V_low
+ 9.615010000e-07 V_low
+ 9.616000000e-07 V_low
+ 9.616010000e-07 V_low
+ 9.617000000e-07 V_low
+ 9.617010000e-07 V_low
+ 9.618000000e-07 V_low
+ 9.618010000e-07 V_low
+ 9.619000000e-07 V_low
+ 9.619010000e-07 V_low
+ 9.620000000e-07 V_low
+ 9.620010000e-07 V_low
+ 9.621000000e-07 V_low
+ 9.621010000e-07 V_low
+ 9.622000000e-07 V_low
+ 9.622010000e-07 V_low
+ 9.623000000e-07 V_low
+ 9.623010000e-07 V_low
+ 9.624000000e-07 V_low
+ 9.624010000e-07 V_low
+ 9.625000000e-07 V_low
+ 9.625010000e-07 V_low
+ 9.626000000e-07 V_low
+ 9.626010000e-07 V_low
+ 9.627000000e-07 V_low
+ 9.627010000e-07 V_low
+ 9.628000000e-07 V_low
+ 9.628010000e-07 V_low
+ 9.629000000e-07 V_low
+ 9.629010000e-07 V_low
+ 9.630000000e-07 V_low
+ 9.630010000e-07 V_low
+ 9.631000000e-07 V_low
+ 9.631010000e-07 V_low
+ 9.632000000e-07 V_low
+ 9.632010000e-07 V_low
+ 9.633000000e-07 V_low
+ 9.633010000e-07 V_low
+ 9.634000000e-07 V_low
+ 9.634010000e-07 V_low
+ 9.635000000e-07 V_low
+ 9.635010000e-07 V_low
+ 9.636000000e-07 V_low
+ 9.636010000e-07 V_low
+ 9.637000000e-07 V_low
+ 9.637010000e-07 V_low
+ 9.638000000e-07 V_low
+ 9.638010000e-07 V_low
+ 9.639000000e-07 V_low
+ 9.639010000e-07 V_low
+ 9.640000000e-07 V_low
+ 9.640010000e-07 V_low
+ 9.641000000e-07 V_low
+ 9.641010000e-07 V_low
+ 9.642000000e-07 V_low
+ 9.642010000e-07 V_low
+ 9.643000000e-07 V_low
+ 9.643010000e-07 V_low
+ 9.644000000e-07 V_low
+ 9.644010000e-07 V_low
+ 9.645000000e-07 V_low
+ 9.645010000e-07 V_low
+ 9.646000000e-07 V_low
+ 9.646010000e-07 V_low
+ 9.647000000e-07 V_low
+ 9.647010000e-07 V_low
+ 9.648000000e-07 V_low
+ 9.648010000e-07 V_low
+ 9.649000000e-07 V_low
+ 9.649010000e-07 V_hig
+ 9.650000000e-07 V_hig
+ 9.650010000e-07 V_hig
+ 9.651000000e-07 V_hig
+ 9.651010000e-07 V_hig
+ 9.652000000e-07 V_hig
+ 9.652010000e-07 V_hig
+ 9.653000000e-07 V_hig
+ 9.653010000e-07 V_hig
+ 9.654000000e-07 V_hig
+ 9.654010000e-07 V_hig
+ 9.655000000e-07 V_hig
+ 9.655010000e-07 V_hig
+ 9.656000000e-07 V_hig
+ 9.656010000e-07 V_hig
+ 9.657000000e-07 V_hig
+ 9.657010000e-07 V_hig
+ 9.658000000e-07 V_hig
+ 9.658010000e-07 V_hig
+ 9.659000000e-07 V_hig
+ 9.659010000e-07 V_hig
+ 9.660000000e-07 V_hig
+ 9.660010000e-07 V_hig
+ 9.661000000e-07 V_hig
+ 9.661010000e-07 V_hig
+ 9.662000000e-07 V_hig
+ 9.662010000e-07 V_hig
+ 9.663000000e-07 V_hig
+ 9.663010000e-07 V_hig
+ 9.664000000e-07 V_hig
+ 9.664010000e-07 V_hig
+ 9.665000000e-07 V_hig
+ 9.665010000e-07 V_hig
+ 9.666000000e-07 V_hig
+ 9.666010000e-07 V_hig
+ 9.667000000e-07 V_hig
+ 9.667010000e-07 V_hig
+ 9.668000000e-07 V_hig
+ 9.668010000e-07 V_hig
+ 9.669000000e-07 V_hig
+ 9.669010000e-07 V_hig
+ 9.670000000e-07 V_hig
+ 9.670010000e-07 V_hig
+ 9.671000000e-07 V_hig
+ 9.671010000e-07 V_hig
+ 9.672000000e-07 V_hig
+ 9.672010000e-07 V_hig
+ 9.673000000e-07 V_hig
+ 9.673010000e-07 V_hig
+ 9.674000000e-07 V_hig
+ 9.674010000e-07 V_hig
+ 9.675000000e-07 V_hig
+ 9.675010000e-07 V_hig
+ 9.676000000e-07 V_hig
+ 9.676010000e-07 V_hig
+ 9.677000000e-07 V_hig
+ 9.677010000e-07 V_hig
+ 9.678000000e-07 V_hig
+ 9.678010000e-07 V_hig
+ 9.679000000e-07 V_hig
+ 9.679010000e-07 V_hig
+ 9.680000000e-07 V_hig
+ 9.680010000e-07 V_hig
+ 9.681000000e-07 V_hig
+ 9.681010000e-07 V_hig
+ 9.682000000e-07 V_hig
+ 9.682010000e-07 V_hig
+ 9.683000000e-07 V_hig
+ 9.683010000e-07 V_hig
+ 9.684000000e-07 V_hig
+ 9.684010000e-07 V_hig
+ 9.685000000e-07 V_hig
+ 9.685010000e-07 V_hig
+ 9.686000000e-07 V_hig
+ 9.686010000e-07 V_hig
+ 9.687000000e-07 V_hig
+ 9.687010000e-07 V_hig
+ 9.688000000e-07 V_hig
+ 9.688010000e-07 V_hig
+ 9.689000000e-07 V_hig
+ 9.689010000e-07 V_low
+ 9.690000000e-07 V_low
+ 9.690010000e-07 V_low
+ 9.691000000e-07 V_low
+ 9.691010000e-07 V_low
+ 9.692000000e-07 V_low
+ 9.692010000e-07 V_low
+ 9.693000000e-07 V_low
+ 9.693010000e-07 V_low
+ 9.694000000e-07 V_low
+ 9.694010000e-07 V_low
+ 9.695000000e-07 V_low
+ 9.695010000e-07 V_low
+ 9.696000000e-07 V_low
+ 9.696010000e-07 V_low
+ 9.697000000e-07 V_low
+ 9.697010000e-07 V_low
+ 9.698000000e-07 V_low
+ 9.698010000e-07 V_low
+ 9.699000000e-07 V_low
+ 9.699010000e-07 V_low
+ 9.700000000e-07 V_low
+ 9.700010000e-07 V_low
+ 9.701000000e-07 V_low
+ 9.701010000e-07 V_low
+ 9.702000000e-07 V_low
+ 9.702010000e-07 V_low
+ 9.703000000e-07 V_low
+ 9.703010000e-07 V_low
+ 9.704000000e-07 V_low
+ 9.704010000e-07 V_low
+ 9.705000000e-07 V_low
+ 9.705010000e-07 V_low
+ 9.706000000e-07 V_low
+ 9.706010000e-07 V_low
+ 9.707000000e-07 V_low
+ 9.707010000e-07 V_low
+ 9.708000000e-07 V_low
+ 9.708010000e-07 V_low
+ 9.709000000e-07 V_low
+ 9.709010000e-07 V_hig
+ 9.710000000e-07 V_hig
+ 9.710010000e-07 V_hig
+ 9.711000000e-07 V_hig
+ 9.711010000e-07 V_hig
+ 9.712000000e-07 V_hig
+ 9.712010000e-07 V_hig
+ 9.713000000e-07 V_hig
+ 9.713010000e-07 V_hig
+ 9.714000000e-07 V_hig
+ 9.714010000e-07 V_hig
+ 9.715000000e-07 V_hig
+ 9.715010000e-07 V_hig
+ 9.716000000e-07 V_hig
+ 9.716010000e-07 V_hig
+ 9.717000000e-07 V_hig
+ 9.717010000e-07 V_hig
+ 9.718000000e-07 V_hig
+ 9.718010000e-07 V_hig
+ 9.719000000e-07 V_hig
+ 9.719010000e-07 V_low
+ 9.720000000e-07 V_low
+ 9.720010000e-07 V_low
+ 9.721000000e-07 V_low
+ 9.721010000e-07 V_low
+ 9.722000000e-07 V_low
+ 9.722010000e-07 V_low
+ 9.723000000e-07 V_low
+ 9.723010000e-07 V_low
+ 9.724000000e-07 V_low
+ 9.724010000e-07 V_low
+ 9.725000000e-07 V_low
+ 9.725010000e-07 V_low
+ 9.726000000e-07 V_low
+ 9.726010000e-07 V_low
+ 9.727000000e-07 V_low
+ 9.727010000e-07 V_low
+ 9.728000000e-07 V_low
+ 9.728010000e-07 V_low
+ 9.729000000e-07 V_low
+ 9.729010000e-07 V_low
+ 9.730000000e-07 V_low
+ 9.730010000e-07 V_low
+ 9.731000000e-07 V_low
+ 9.731010000e-07 V_low
+ 9.732000000e-07 V_low
+ 9.732010000e-07 V_low
+ 9.733000000e-07 V_low
+ 9.733010000e-07 V_low
+ 9.734000000e-07 V_low
+ 9.734010000e-07 V_low
+ 9.735000000e-07 V_low
+ 9.735010000e-07 V_low
+ 9.736000000e-07 V_low
+ 9.736010000e-07 V_low
+ 9.737000000e-07 V_low
+ 9.737010000e-07 V_low
+ 9.738000000e-07 V_low
+ 9.738010000e-07 V_low
+ 9.739000000e-07 V_low
+ 9.739010000e-07 V_low
+ 9.740000000e-07 V_low
+ 9.740010000e-07 V_low
+ 9.741000000e-07 V_low
+ 9.741010000e-07 V_low
+ 9.742000000e-07 V_low
+ 9.742010000e-07 V_low
+ 9.743000000e-07 V_low
+ 9.743010000e-07 V_low
+ 9.744000000e-07 V_low
+ 9.744010000e-07 V_low
+ 9.745000000e-07 V_low
+ 9.745010000e-07 V_low
+ 9.746000000e-07 V_low
+ 9.746010000e-07 V_low
+ 9.747000000e-07 V_low
+ 9.747010000e-07 V_low
+ 9.748000000e-07 V_low
+ 9.748010000e-07 V_low
+ 9.749000000e-07 V_low
+ 9.749010000e-07 V_hig
+ 9.750000000e-07 V_hig
+ 9.750010000e-07 V_hig
+ 9.751000000e-07 V_hig
+ 9.751010000e-07 V_hig
+ 9.752000000e-07 V_hig
+ 9.752010000e-07 V_hig
+ 9.753000000e-07 V_hig
+ 9.753010000e-07 V_hig
+ 9.754000000e-07 V_hig
+ 9.754010000e-07 V_hig
+ 9.755000000e-07 V_hig
+ 9.755010000e-07 V_hig
+ 9.756000000e-07 V_hig
+ 9.756010000e-07 V_hig
+ 9.757000000e-07 V_hig
+ 9.757010000e-07 V_hig
+ 9.758000000e-07 V_hig
+ 9.758010000e-07 V_hig
+ 9.759000000e-07 V_hig
+ 9.759010000e-07 V_hig
+ 9.760000000e-07 V_hig
+ 9.760010000e-07 V_hig
+ 9.761000000e-07 V_hig
+ 9.761010000e-07 V_hig
+ 9.762000000e-07 V_hig
+ 9.762010000e-07 V_hig
+ 9.763000000e-07 V_hig
+ 9.763010000e-07 V_hig
+ 9.764000000e-07 V_hig
+ 9.764010000e-07 V_hig
+ 9.765000000e-07 V_hig
+ 9.765010000e-07 V_hig
+ 9.766000000e-07 V_hig
+ 9.766010000e-07 V_hig
+ 9.767000000e-07 V_hig
+ 9.767010000e-07 V_hig
+ 9.768000000e-07 V_hig
+ 9.768010000e-07 V_hig
+ 9.769000000e-07 V_hig
+ 9.769010000e-07 V_low
+ 9.770000000e-07 V_low
+ 9.770010000e-07 V_low
+ 9.771000000e-07 V_low
+ 9.771010000e-07 V_low
+ 9.772000000e-07 V_low
+ 9.772010000e-07 V_low
+ 9.773000000e-07 V_low
+ 9.773010000e-07 V_low
+ 9.774000000e-07 V_low
+ 9.774010000e-07 V_low
+ 9.775000000e-07 V_low
+ 9.775010000e-07 V_low
+ 9.776000000e-07 V_low
+ 9.776010000e-07 V_low
+ 9.777000000e-07 V_low
+ 9.777010000e-07 V_low
+ 9.778000000e-07 V_low
+ 9.778010000e-07 V_low
+ 9.779000000e-07 V_low
+ 9.779010000e-07 V_hig
+ 9.780000000e-07 V_hig
+ 9.780010000e-07 V_hig
+ 9.781000000e-07 V_hig
+ 9.781010000e-07 V_hig
+ 9.782000000e-07 V_hig
+ 9.782010000e-07 V_hig
+ 9.783000000e-07 V_hig
+ 9.783010000e-07 V_hig
+ 9.784000000e-07 V_hig
+ 9.784010000e-07 V_hig
+ 9.785000000e-07 V_hig
+ 9.785010000e-07 V_hig
+ 9.786000000e-07 V_hig
+ 9.786010000e-07 V_hig
+ 9.787000000e-07 V_hig
+ 9.787010000e-07 V_hig
+ 9.788000000e-07 V_hig
+ 9.788010000e-07 V_hig
+ 9.789000000e-07 V_hig
+ 9.789010000e-07 V_hig
+ 9.790000000e-07 V_hig
+ 9.790010000e-07 V_hig
+ 9.791000000e-07 V_hig
+ 9.791010000e-07 V_hig
+ 9.792000000e-07 V_hig
+ 9.792010000e-07 V_hig
+ 9.793000000e-07 V_hig
+ 9.793010000e-07 V_hig
+ 9.794000000e-07 V_hig
+ 9.794010000e-07 V_hig
+ 9.795000000e-07 V_hig
+ 9.795010000e-07 V_hig
+ 9.796000000e-07 V_hig
+ 9.796010000e-07 V_hig
+ 9.797000000e-07 V_hig
+ 9.797010000e-07 V_hig
+ 9.798000000e-07 V_hig
+ 9.798010000e-07 V_hig
+ 9.799000000e-07 V_hig
+ 9.799010000e-07 V_low
+ 9.800000000e-07 V_low
+ 9.800010000e-07 V_low
+ 9.801000000e-07 V_low
+ 9.801010000e-07 V_low
+ 9.802000000e-07 V_low
+ 9.802010000e-07 V_low
+ 9.803000000e-07 V_low
+ 9.803010000e-07 V_low
+ 9.804000000e-07 V_low
+ 9.804010000e-07 V_low
+ 9.805000000e-07 V_low
+ 9.805010000e-07 V_low
+ 9.806000000e-07 V_low
+ 9.806010000e-07 V_low
+ 9.807000000e-07 V_low
+ 9.807010000e-07 V_low
+ 9.808000000e-07 V_low
+ 9.808010000e-07 V_low
+ 9.809000000e-07 V_low
+ 9.809010000e-07 V_low
+ 9.810000000e-07 V_low
+ 9.810010000e-07 V_low
+ 9.811000000e-07 V_low
+ 9.811010000e-07 V_low
+ 9.812000000e-07 V_low
+ 9.812010000e-07 V_low
+ 9.813000000e-07 V_low
+ 9.813010000e-07 V_low
+ 9.814000000e-07 V_low
+ 9.814010000e-07 V_low
+ 9.815000000e-07 V_low
+ 9.815010000e-07 V_low
+ 9.816000000e-07 V_low
+ 9.816010000e-07 V_low
+ 9.817000000e-07 V_low
+ 9.817010000e-07 V_low
+ 9.818000000e-07 V_low
+ 9.818010000e-07 V_low
+ 9.819000000e-07 V_low
+ 9.819010000e-07 V_hig
+ 9.820000000e-07 V_hig
+ 9.820010000e-07 V_hig
+ 9.821000000e-07 V_hig
+ 9.821010000e-07 V_hig
+ 9.822000000e-07 V_hig
+ 9.822010000e-07 V_hig
+ 9.823000000e-07 V_hig
+ 9.823010000e-07 V_hig
+ 9.824000000e-07 V_hig
+ 9.824010000e-07 V_hig
+ 9.825000000e-07 V_hig
+ 9.825010000e-07 V_hig
+ 9.826000000e-07 V_hig
+ 9.826010000e-07 V_hig
+ 9.827000000e-07 V_hig
+ 9.827010000e-07 V_hig
+ 9.828000000e-07 V_hig
+ 9.828010000e-07 V_hig
+ 9.829000000e-07 V_hig
+ 9.829010000e-07 V_low
+ 9.830000000e-07 V_low
+ 9.830010000e-07 V_low
+ 9.831000000e-07 V_low
+ 9.831010000e-07 V_low
+ 9.832000000e-07 V_low
+ 9.832010000e-07 V_low
+ 9.833000000e-07 V_low
+ 9.833010000e-07 V_low
+ 9.834000000e-07 V_low
+ 9.834010000e-07 V_low
+ 9.835000000e-07 V_low
+ 9.835010000e-07 V_low
+ 9.836000000e-07 V_low
+ 9.836010000e-07 V_low
+ 9.837000000e-07 V_low
+ 9.837010000e-07 V_low
+ 9.838000000e-07 V_low
+ 9.838010000e-07 V_low
+ 9.839000000e-07 V_low
+ 9.839010000e-07 V_low
+ 9.840000000e-07 V_low
+ 9.840010000e-07 V_low
+ 9.841000000e-07 V_low
+ 9.841010000e-07 V_low
+ 9.842000000e-07 V_low
+ 9.842010000e-07 V_low
+ 9.843000000e-07 V_low
+ 9.843010000e-07 V_low
+ 9.844000000e-07 V_low
+ 9.844010000e-07 V_low
+ 9.845000000e-07 V_low
+ 9.845010000e-07 V_low
+ 9.846000000e-07 V_low
+ 9.846010000e-07 V_low
+ 9.847000000e-07 V_low
+ 9.847010000e-07 V_low
+ 9.848000000e-07 V_low
+ 9.848010000e-07 V_low
+ 9.849000000e-07 V_low
+ 9.849010000e-07 V_low
+ 9.850000000e-07 V_low
+ 9.850010000e-07 V_low
+ 9.851000000e-07 V_low
+ 9.851010000e-07 V_low
+ 9.852000000e-07 V_low
+ 9.852010000e-07 V_low
+ 9.853000000e-07 V_low
+ 9.853010000e-07 V_low
+ 9.854000000e-07 V_low
+ 9.854010000e-07 V_low
+ 9.855000000e-07 V_low
+ 9.855010000e-07 V_low
+ 9.856000000e-07 V_low
+ 9.856010000e-07 V_low
+ 9.857000000e-07 V_low
+ 9.857010000e-07 V_low
+ 9.858000000e-07 V_low
+ 9.858010000e-07 V_low
+ 9.859000000e-07 V_low
+ 9.859010000e-07 V_hig
+ 9.860000000e-07 V_hig
+ 9.860010000e-07 V_hig
+ 9.861000000e-07 V_hig
+ 9.861010000e-07 V_hig
+ 9.862000000e-07 V_hig
+ 9.862010000e-07 V_hig
+ 9.863000000e-07 V_hig
+ 9.863010000e-07 V_hig
+ 9.864000000e-07 V_hig
+ 9.864010000e-07 V_hig
+ 9.865000000e-07 V_hig
+ 9.865010000e-07 V_hig
+ 9.866000000e-07 V_hig
+ 9.866010000e-07 V_hig
+ 9.867000000e-07 V_hig
+ 9.867010000e-07 V_hig
+ 9.868000000e-07 V_hig
+ 9.868010000e-07 V_hig
+ 9.869000000e-07 V_hig
+ 9.869010000e-07 V_hig
+ 9.870000000e-07 V_hig
+ 9.870010000e-07 V_hig
+ 9.871000000e-07 V_hig
+ 9.871010000e-07 V_hig
+ 9.872000000e-07 V_hig
+ 9.872010000e-07 V_hig
+ 9.873000000e-07 V_hig
+ 9.873010000e-07 V_hig
+ 9.874000000e-07 V_hig
+ 9.874010000e-07 V_hig
+ 9.875000000e-07 V_hig
+ 9.875010000e-07 V_hig
+ 9.876000000e-07 V_hig
+ 9.876010000e-07 V_hig
+ 9.877000000e-07 V_hig
+ 9.877010000e-07 V_hig
+ 9.878000000e-07 V_hig
+ 9.878010000e-07 V_hig
+ 9.879000000e-07 V_hig
+ 9.879010000e-07 V_low
+ 9.880000000e-07 V_low
+ 9.880010000e-07 V_low
+ 9.881000000e-07 V_low
+ 9.881010000e-07 V_low
+ 9.882000000e-07 V_low
+ 9.882010000e-07 V_low
+ 9.883000000e-07 V_low
+ 9.883010000e-07 V_low
+ 9.884000000e-07 V_low
+ 9.884010000e-07 V_low
+ 9.885000000e-07 V_low
+ 9.885010000e-07 V_low
+ 9.886000000e-07 V_low
+ 9.886010000e-07 V_low
+ 9.887000000e-07 V_low
+ 9.887010000e-07 V_low
+ 9.888000000e-07 V_low
+ 9.888010000e-07 V_low
+ 9.889000000e-07 V_low
+ 9.889010000e-07 V_hig
+ 9.890000000e-07 V_hig
+ 9.890010000e-07 V_hig
+ 9.891000000e-07 V_hig
+ 9.891010000e-07 V_hig
+ 9.892000000e-07 V_hig
+ 9.892010000e-07 V_hig
+ 9.893000000e-07 V_hig
+ 9.893010000e-07 V_hig
+ 9.894000000e-07 V_hig
+ 9.894010000e-07 V_hig
+ 9.895000000e-07 V_hig
+ 9.895010000e-07 V_hig
+ 9.896000000e-07 V_hig
+ 9.896010000e-07 V_hig
+ 9.897000000e-07 V_hig
+ 9.897010000e-07 V_hig
+ 9.898000000e-07 V_hig
+ 9.898010000e-07 V_hig
+ 9.899000000e-07 V_hig
+ 9.899010000e-07 V_hig
+ 9.900000000e-07 V_hig
+ 9.900010000e-07 V_hig
+ 9.901000000e-07 V_hig
+ 9.901010000e-07 V_hig
+ 9.902000000e-07 V_hig
+ 9.902010000e-07 V_hig
+ 9.903000000e-07 V_hig
+ 9.903010000e-07 V_hig
+ 9.904000000e-07 V_hig
+ 9.904010000e-07 V_hig
+ 9.905000000e-07 V_hig
+ 9.905010000e-07 V_hig
+ 9.906000000e-07 V_hig
+ 9.906010000e-07 V_hig
+ 9.907000000e-07 V_hig
+ 9.907010000e-07 V_hig
+ 9.908000000e-07 V_hig
+ 9.908010000e-07 V_hig
+ 9.909000000e-07 V_hig
+ 9.909010000e-07 V_hig
+ 9.910000000e-07 V_hig
+ 9.910010000e-07 V_hig
+ 9.911000000e-07 V_hig
+ 9.911010000e-07 V_hig
+ 9.912000000e-07 V_hig
+ 9.912010000e-07 V_hig
+ 9.913000000e-07 V_hig
+ 9.913010000e-07 V_hig
+ 9.914000000e-07 V_hig
+ 9.914010000e-07 V_hig
+ 9.915000000e-07 V_hig
+ 9.915010000e-07 V_hig
+ 9.916000000e-07 V_hig
+ 9.916010000e-07 V_hig
+ 9.917000000e-07 V_hig
+ 9.917010000e-07 V_hig
+ 9.918000000e-07 V_hig
+ 9.918010000e-07 V_hig
+ 9.919000000e-07 V_hig
+ 9.919010000e-07 V_low
+ 9.920000000e-07 V_low
+ 9.920010000e-07 V_low
+ 9.921000000e-07 V_low
+ 9.921010000e-07 V_low
+ 9.922000000e-07 V_low
+ 9.922010000e-07 V_low
+ 9.923000000e-07 V_low
+ 9.923010000e-07 V_low
+ 9.924000000e-07 V_low
+ 9.924010000e-07 V_low
+ 9.925000000e-07 V_low
+ 9.925010000e-07 V_low
+ 9.926000000e-07 V_low
+ 9.926010000e-07 V_low
+ 9.927000000e-07 V_low
+ 9.927010000e-07 V_low
+ 9.928000000e-07 V_low
+ 9.928010000e-07 V_low
+ 9.929000000e-07 V_low
+ 9.929010000e-07 V_hig
+ 9.930000000e-07 V_hig
+ 9.930010000e-07 V_hig
+ 9.931000000e-07 V_hig
+ 9.931010000e-07 V_hig
+ 9.932000000e-07 V_hig
+ 9.932010000e-07 V_hig
+ 9.933000000e-07 V_hig
+ 9.933010000e-07 V_hig
+ 9.934000000e-07 V_hig
+ 9.934010000e-07 V_hig
+ 9.935000000e-07 V_hig
+ 9.935010000e-07 V_hig
+ 9.936000000e-07 V_hig
+ 9.936010000e-07 V_hig
+ 9.937000000e-07 V_hig
+ 9.937010000e-07 V_hig
+ 9.938000000e-07 V_hig
+ 9.938010000e-07 V_hig
+ 9.939000000e-07 V_hig
+ 9.939010000e-07 V_low
+ 9.940000000e-07 V_low
+ 9.940010000e-07 V_low
+ 9.941000000e-07 V_low
+ 9.941010000e-07 V_low
+ 9.942000000e-07 V_low
+ 9.942010000e-07 V_low
+ 9.943000000e-07 V_low
+ 9.943010000e-07 V_low
+ 9.944000000e-07 V_low
+ 9.944010000e-07 V_low
+ 9.945000000e-07 V_low
+ 9.945010000e-07 V_low
+ 9.946000000e-07 V_low
+ 9.946010000e-07 V_low
+ 9.947000000e-07 V_low
+ 9.947010000e-07 V_low
+ 9.948000000e-07 V_low
+ 9.948010000e-07 V_low
+ 9.949000000e-07 V_low
+ 9.949010000e-07 V_hig
+ 9.950000000e-07 V_hig
+ 9.950010000e-07 V_hig
+ 9.951000000e-07 V_hig
+ 9.951010000e-07 V_hig
+ 9.952000000e-07 V_hig
+ 9.952010000e-07 V_hig
+ 9.953000000e-07 V_hig
+ 9.953010000e-07 V_hig
+ 9.954000000e-07 V_hig
+ 9.954010000e-07 V_hig
+ 9.955000000e-07 V_hig
+ 9.955010000e-07 V_hig
+ 9.956000000e-07 V_hig
+ 9.956010000e-07 V_hig
+ 9.957000000e-07 V_hig
+ 9.957010000e-07 V_hig
+ 9.958000000e-07 V_hig
+ 9.958010000e-07 V_hig
+ 9.959000000e-07 V_hig
+ 9.959010000e-07 V_low
+ 9.960000000e-07 V_low
+ 9.960010000e-07 V_low
+ 9.961000000e-07 V_low
+ 9.961010000e-07 V_low
+ 9.962000000e-07 V_low
+ 9.962010000e-07 V_low
+ 9.963000000e-07 V_low
+ 9.963010000e-07 V_low
+ 9.964000000e-07 V_low
+ 9.964010000e-07 V_low
+ 9.965000000e-07 V_low
+ 9.965010000e-07 V_low
+ 9.966000000e-07 V_low
+ 9.966010000e-07 V_low
+ 9.967000000e-07 V_low
+ 9.967010000e-07 V_low
+ 9.968000000e-07 V_low
+ 9.968010000e-07 V_low
+ 9.969000000e-07 V_low
+ 9.969010000e-07 V_low
+ 9.970000000e-07 V_low
+ 9.970010000e-07 V_low
+ 9.971000000e-07 V_low
+ 9.971010000e-07 V_low
+ 9.972000000e-07 V_low
+ 9.972010000e-07 V_low
+ 9.973000000e-07 V_low
+ 9.973010000e-07 V_low
+ 9.974000000e-07 V_low
+ 9.974010000e-07 V_low
+ 9.975000000e-07 V_low
+ 9.975010000e-07 V_low
+ 9.976000000e-07 V_low
+ 9.976010000e-07 V_low
+ 9.977000000e-07 V_low
+ 9.977010000e-07 V_low
+ 9.978000000e-07 V_low
+ 9.978010000e-07 V_low
+ 9.979000000e-07 V_low
+ 9.979010000e-07 V_hig
+ 9.980000000e-07 V_hig
+ 9.980010000e-07 V_hig
+ 9.981000000e-07 V_hig
+ 9.981010000e-07 V_hig
+ 9.982000000e-07 V_hig
+ 9.982010000e-07 V_hig
+ 9.983000000e-07 V_hig
+ 9.983010000e-07 V_hig
+ 9.984000000e-07 V_hig
+ 9.984010000e-07 V_hig
+ 9.985000000e-07 V_hig
+ 9.985010000e-07 V_hig
+ 9.986000000e-07 V_hig
+ 9.986010000e-07 V_hig
+ 9.987000000e-07 V_hig
+ 9.987010000e-07 V_hig
+ 9.988000000e-07 V_hig
+ 9.988010000e-07 V_hig
+ 9.989000000e-07 V_hig
+ 9.989010000e-07 V_low
+ 9.990000000e-07 V_low
+ 9.990010000e-07 V_low
+ 9.991000000e-07 V_low
+ 9.991010000e-07 V_low
+ 9.992000000e-07 V_low
+ 9.992010000e-07 V_low
+ 9.993000000e-07 V_low
+ 9.993010000e-07 V_low
+ 9.994000000e-07 V_low
+ 9.994010000e-07 V_low
+ 9.995000000e-07 V_low
+ 9.995010000e-07 V_low
+ 9.996000000e-07 V_low
+ 9.996010000e-07 V_low
+ 9.997000000e-07 V_low
+ 9.997010000e-07 V_low
+ 9.998000000e-07 V_low
+ 9.998010000e-07 V_low
+ 9.999000000e-07 V_low
+ 9.999010000e-07 V_low
+ 1.000000000e-06 V_low
+ 1.000001000e-06 V_low
+ 1.000100000e-06 V_low
+ 1.000101000e-06 V_low
+ 1.000200000e-06 V_low
+ 1.000201000e-06 V_low
+ 1.000300000e-06 V_low
+ 1.000301000e-06 V_low
+ 1.000400000e-06 V_low
+ 1.000401000e-06 V_low
+ 1.000500000e-06 V_low
+ 1.000501000e-06 V_low
+ 1.000600000e-06 V_low
+ 1.000601000e-06 V_low
+ 1.000700000e-06 V_low
+ 1.000701000e-06 V_low
+ 1.000800000e-06 V_low
+ 1.000801000e-06 V_low
+ 1.000900000e-06 V_low
+ 
v1 a 0 PWL
+ 1.000000000e-12 V_low
+ 1.000000000e-09 V_low
+ 1.001000000e-09 V_low
+ 1.100000000e-09 V_low
+ 1.101000000e-09 V_low
+ 1.200000000e-09 V_low
+ 1.201000000e-09 V_low
+ 1.300000000e-09 V_low
+ 1.301000000e-09 V_low
+ 1.400000000e-09 V_low
+ 1.401000000e-09 V_low
+ 1.500000000e-09 V_low
+ 1.501000000e-09 V_low
+ 1.600000000e-09 V_low
+ 1.601000000e-09 V_low
+ 1.700000000e-09 V_low
+ 1.701000000e-09 V_low
+ 1.800000000e-09 V_low
+ 1.801000000e-09 V_low
+ 1.900000000e-09 V_low
+ 1.901000000e-09 V_hig
+ 2.000000000e-09 V_hig
+ 2.001000000e-09 V_hig
+ 2.100000000e-09 V_hig
+ 2.101000000e-09 V_hig
+ 2.200000000e-09 V_hig
+ 2.201000000e-09 V_hig
+ 2.300000000e-09 V_hig
+ 2.301000000e-09 V_hig
+ 2.400000000e-09 V_hig
+ 2.401000000e-09 V_hig
+ 2.500000000e-09 V_hig
+ 2.501000000e-09 V_hig
+ 2.600000000e-09 V_hig
+ 2.601000000e-09 V_hig
+ 2.700000000e-09 V_hig
+ 2.701000000e-09 V_hig
+ 2.800000000e-09 V_hig
+ 2.801000000e-09 V_hig
+ 2.900000000e-09 V_hig
+ 2.901000000e-09 V_low
+ 3.000000000e-09 V_low
+ 3.001000000e-09 V_low
+ 3.100000000e-09 V_low
+ 3.101000000e-09 V_low
+ 3.200000000e-09 V_low
+ 3.201000000e-09 V_low
+ 3.300000000e-09 V_low
+ 3.301000000e-09 V_low
+ 3.400000000e-09 V_low
+ 3.401000000e-09 V_low
+ 3.500000000e-09 V_low
+ 3.501000000e-09 V_low
+ 3.600000000e-09 V_low
+ 3.601000000e-09 V_low
+ 3.700000000e-09 V_low
+ 3.701000000e-09 V_low
+ 3.800000000e-09 V_low
+ 3.801000000e-09 V_low
+ 3.900000000e-09 V_low
+ 3.901000000e-09 V_hig
+ 4.000000000e-09 V_hig
+ 4.001000000e-09 V_hig
+ 4.100000000e-09 V_hig
+ 4.101000000e-09 V_hig
+ 4.200000000e-09 V_hig
+ 4.201000000e-09 V_hig
+ 4.300000000e-09 V_hig
+ 4.301000000e-09 V_hig
+ 4.400000000e-09 V_hig
+ 4.401000000e-09 V_hig
+ 4.500000000e-09 V_hig
+ 4.501000000e-09 V_hig
+ 4.600000000e-09 V_hig
+ 4.601000000e-09 V_hig
+ 4.700000000e-09 V_hig
+ 4.701000000e-09 V_hig
+ 4.800000000e-09 V_hig
+ 4.801000000e-09 V_hig
+ 4.900000000e-09 V_hig
+ 4.901000000e-09 V_hig
+ 5.000000000e-09 V_hig
+ 5.001000000e-09 V_hig
+ 5.100000000e-09 V_hig
+ 5.101000000e-09 V_hig
+ 5.200000000e-09 V_hig
+ 5.201000000e-09 V_hig
+ 5.300000000e-09 V_hig
+ 5.301000000e-09 V_hig
+ 5.400000000e-09 V_hig
+ 5.401000000e-09 V_hig
+ 5.500000000e-09 V_hig
+ 5.501000000e-09 V_hig
+ 5.600000000e-09 V_hig
+ 5.601000000e-09 V_hig
+ 5.700000000e-09 V_hig
+ 5.701000000e-09 V_hig
+ 5.800000000e-09 V_hig
+ 5.801000000e-09 V_hig
+ 5.900000000e-09 V_hig
+ 5.901000000e-09 V_low
+ 6.000000000e-09 V_low
+ 6.001000000e-09 V_low
+ 6.100000000e-09 V_low
+ 6.101000000e-09 V_low
+ 6.200000000e-09 V_low
+ 6.201000000e-09 V_low
+ 6.300000000e-09 V_low
+ 6.301000000e-09 V_low
+ 6.400000000e-09 V_low
+ 6.401000000e-09 V_low
+ 6.500000000e-09 V_low
+ 6.501000000e-09 V_low
+ 6.600000000e-09 V_low
+ 6.601000000e-09 V_low
+ 6.700000000e-09 V_low
+ 6.701000000e-09 V_low
+ 6.800000000e-09 V_low
+ 6.801000000e-09 V_low
+ 6.900000000e-09 V_low
+ 6.901000000e-09 V_low
+ 7.000000000e-09 V_low
+ 7.001000000e-09 V_low
+ 7.100000000e-09 V_low
+ 7.101000000e-09 V_low
+ 7.200000000e-09 V_low
+ 7.201000000e-09 V_low
+ 7.300000000e-09 V_low
+ 7.301000000e-09 V_low
+ 7.400000000e-09 V_low
+ 7.401000000e-09 V_low
+ 7.500000000e-09 V_low
+ 7.501000000e-09 V_low
+ 7.600000000e-09 V_low
+ 7.601000000e-09 V_low
+ 7.700000000e-09 V_low
+ 7.701000000e-09 V_low
+ 7.800000000e-09 V_low
+ 7.801000000e-09 V_low
+ 7.900000000e-09 V_low
+ 7.901000000e-09 V_hig
+ 8.000000000e-09 V_hig
+ 8.001000000e-09 V_hig
+ 8.100000000e-09 V_hig
+ 8.101000000e-09 V_hig
+ 8.200000000e-09 V_hig
+ 8.201000000e-09 V_hig
+ 8.300000000e-09 V_hig
+ 8.301000000e-09 V_hig
+ 8.400000000e-09 V_hig
+ 8.401000000e-09 V_hig
+ 8.500000000e-09 V_hig
+ 8.501000000e-09 V_hig
+ 8.600000000e-09 V_hig
+ 8.601000000e-09 V_hig
+ 8.700000000e-09 V_hig
+ 8.701000000e-09 V_hig
+ 8.800000000e-09 V_hig
+ 8.801000000e-09 V_hig
+ 8.900000000e-09 V_hig
+ 8.901000000e-09 V_low
+ 9.000000000e-09 V_low
+ 9.001000000e-09 V_low
+ 9.100000000e-09 V_low
+ 9.101000000e-09 V_low
+ 9.200000000e-09 V_low
+ 9.201000000e-09 V_low
+ 9.300000000e-09 V_low
+ 9.301000000e-09 V_low
+ 9.400000000e-09 V_low
+ 9.401000000e-09 V_low
+ 9.500000000e-09 V_low
+ 9.501000000e-09 V_low
+ 9.600000000e-09 V_low
+ 9.601000000e-09 V_low
+ 9.700000000e-09 V_low
+ 9.701000000e-09 V_low
+ 9.800000000e-09 V_low
+ 9.801000000e-09 V_low
+ 9.900000000e-09 V_low
+ 9.901000000e-09 V_low
+ 1.000000000e-08 V_low
+ 1.000100000e-08 V_low
+ 1.010000000e-08 V_low
+ 1.010100000e-08 V_low
+ 1.020000000e-08 V_low
+ 1.020100000e-08 V_low
+ 1.030000000e-08 V_low
+ 1.030100000e-08 V_low
+ 1.040000000e-08 V_low
+ 1.040100000e-08 V_low
+ 1.050000000e-08 V_low
+ 1.050100000e-08 V_low
+ 1.060000000e-08 V_low
+ 1.060100000e-08 V_low
+ 1.070000000e-08 V_low
+ 1.070100000e-08 V_low
+ 1.080000000e-08 V_low
+ 1.080100000e-08 V_low
+ 1.090000000e-08 V_low
+ 1.090100000e-08 V_hig
+ 1.100000000e-08 V_hig
+ 1.100100000e-08 V_hig
+ 1.110000000e-08 V_hig
+ 1.110100000e-08 V_hig
+ 1.120000000e-08 V_hig
+ 1.120100000e-08 V_hig
+ 1.130000000e-08 V_hig
+ 1.130100000e-08 V_hig
+ 1.140000000e-08 V_hig
+ 1.140100000e-08 V_hig
+ 1.150000000e-08 V_hig
+ 1.150100000e-08 V_hig
+ 1.160000000e-08 V_hig
+ 1.160100000e-08 V_hig
+ 1.170000000e-08 V_hig
+ 1.170100000e-08 V_hig
+ 1.180000000e-08 V_hig
+ 1.180100000e-08 V_hig
+ 1.190000000e-08 V_hig
+ 1.190100000e-08 V_low
+ 1.200000000e-08 V_low
+ 1.200100000e-08 V_low
+ 1.210000000e-08 V_low
+ 1.210100000e-08 V_low
+ 1.220000000e-08 V_low
+ 1.220100000e-08 V_low
+ 1.230000000e-08 V_low
+ 1.230100000e-08 V_low
+ 1.240000000e-08 V_low
+ 1.240100000e-08 V_low
+ 1.250000000e-08 V_low
+ 1.250100000e-08 V_low
+ 1.260000000e-08 V_low
+ 1.260100000e-08 V_low
+ 1.270000000e-08 V_low
+ 1.270100000e-08 V_low
+ 1.280000000e-08 V_low
+ 1.280100000e-08 V_low
+ 1.290000000e-08 V_low
+ 1.290100000e-08 V_hig
+ 1.300000000e-08 V_hig
+ 1.300100000e-08 V_hig
+ 1.310000000e-08 V_hig
+ 1.310100000e-08 V_hig
+ 1.320000000e-08 V_hig
+ 1.320100000e-08 V_hig
+ 1.330000000e-08 V_hig
+ 1.330100000e-08 V_hig
+ 1.340000000e-08 V_hig
+ 1.340100000e-08 V_hig
+ 1.350000000e-08 V_hig
+ 1.350100000e-08 V_hig
+ 1.360000000e-08 V_hig
+ 1.360100000e-08 V_hig
+ 1.370000000e-08 V_hig
+ 1.370100000e-08 V_hig
+ 1.380000000e-08 V_hig
+ 1.380100000e-08 V_hig
+ 1.390000000e-08 V_hig
+ 1.390100000e-08 V_hig
+ 1.400000000e-08 V_hig
+ 1.400100000e-08 V_hig
+ 1.410000000e-08 V_hig
+ 1.410100000e-08 V_hig
+ 1.420000000e-08 V_hig
+ 1.420100000e-08 V_hig
+ 1.430000000e-08 V_hig
+ 1.430100000e-08 V_hig
+ 1.440000000e-08 V_hig
+ 1.440100000e-08 V_hig
+ 1.450000000e-08 V_hig
+ 1.450100000e-08 V_hig
+ 1.460000000e-08 V_hig
+ 1.460100000e-08 V_hig
+ 1.470000000e-08 V_hig
+ 1.470100000e-08 V_hig
+ 1.480000000e-08 V_hig
+ 1.480100000e-08 V_hig
+ 1.490000000e-08 V_hig
+ 1.490100000e-08 V_hig
+ 1.500000000e-08 V_hig
+ 1.500100000e-08 V_hig
+ 1.510000000e-08 V_hig
+ 1.510100000e-08 V_hig
+ 1.520000000e-08 V_hig
+ 1.520100000e-08 V_hig
+ 1.530000000e-08 V_hig
+ 1.530100000e-08 V_hig
+ 1.540000000e-08 V_hig
+ 1.540100000e-08 V_hig
+ 1.550000000e-08 V_hig
+ 1.550100000e-08 V_hig
+ 1.560000000e-08 V_hig
+ 1.560100000e-08 V_hig
+ 1.570000000e-08 V_hig
+ 1.570100000e-08 V_hig
+ 1.580000000e-08 V_hig
+ 1.580100000e-08 V_hig
+ 1.590000000e-08 V_hig
+ 1.590100000e-08 V_hig
+ 1.600000000e-08 V_hig
+ 1.600100000e-08 V_hig
+ 1.610000000e-08 V_hig
+ 1.610100000e-08 V_hig
+ 1.620000000e-08 V_hig
+ 1.620100000e-08 V_hig
+ 1.630000000e-08 V_hig
+ 1.630100000e-08 V_hig
+ 1.640000000e-08 V_hig
+ 1.640100000e-08 V_hig
+ 1.650000000e-08 V_hig
+ 1.650100000e-08 V_hig
+ 1.660000000e-08 V_hig
+ 1.660100000e-08 V_hig
+ 1.670000000e-08 V_hig
+ 1.670100000e-08 V_hig
+ 1.680000000e-08 V_hig
+ 1.680100000e-08 V_hig
+ 1.690000000e-08 V_hig
+ 1.690100000e-08 V_low
+ 1.700000000e-08 V_low
+ 1.700100000e-08 V_low
+ 1.710000000e-08 V_low
+ 1.710100000e-08 V_low
+ 1.720000000e-08 V_low
+ 1.720100000e-08 V_low
+ 1.730000000e-08 V_low
+ 1.730100000e-08 V_low
+ 1.740000000e-08 V_low
+ 1.740100000e-08 V_low
+ 1.750000000e-08 V_low
+ 1.750100000e-08 V_low
+ 1.760000000e-08 V_low
+ 1.760100000e-08 V_low
+ 1.770000000e-08 V_low
+ 1.770100000e-08 V_low
+ 1.780000000e-08 V_low
+ 1.780100000e-08 V_low
+ 1.790000000e-08 V_low
+ 1.790100000e-08 V_hig
+ 1.800000000e-08 V_hig
+ 1.800100000e-08 V_hig
+ 1.810000000e-08 V_hig
+ 1.810100000e-08 V_hig
+ 1.820000000e-08 V_hig
+ 1.820100000e-08 V_hig
+ 1.830000000e-08 V_hig
+ 1.830100000e-08 V_hig
+ 1.840000000e-08 V_hig
+ 1.840100000e-08 V_hig
+ 1.850000000e-08 V_hig
+ 1.850100000e-08 V_hig
+ 1.860000000e-08 V_hig
+ 1.860100000e-08 V_hig
+ 1.870000000e-08 V_hig
+ 1.870100000e-08 V_hig
+ 1.880000000e-08 V_hig
+ 1.880100000e-08 V_hig
+ 1.890000000e-08 V_hig
+ 1.890100000e-08 V_hig
+ 1.900000000e-08 V_hig
+ 1.900100000e-08 V_hig
+ 1.910000000e-08 V_hig
+ 1.910100000e-08 V_hig
+ 1.920000000e-08 V_hig
+ 1.920100000e-08 V_hig
+ 1.930000000e-08 V_hig
+ 1.930100000e-08 V_hig
+ 1.940000000e-08 V_hig
+ 1.940100000e-08 V_hig
+ 1.950000000e-08 V_hig
+ 1.950100000e-08 V_hig
+ 1.960000000e-08 V_hig
+ 1.960100000e-08 V_hig
+ 1.970000000e-08 V_hig
+ 1.970100000e-08 V_hig
+ 1.980000000e-08 V_hig
+ 1.980100000e-08 V_hig
+ 1.990000000e-08 V_hig
+ 1.990100000e-08 V_low
+ 2.000000000e-08 V_low
+ 2.000100000e-08 V_low
+ 2.010000000e-08 V_low
+ 2.010100000e-08 V_low
+ 2.020000000e-08 V_low
+ 2.020100000e-08 V_low
+ 2.030000000e-08 V_low
+ 2.030100000e-08 V_low
+ 2.040000000e-08 V_low
+ 2.040100000e-08 V_low
+ 2.050000000e-08 V_low
+ 2.050100000e-08 V_low
+ 2.060000000e-08 V_low
+ 2.060100000e-08 V_low
+ 2.070000000e-08 V_low
+ 2.070100000e-08 V_low
+ 2.080000000e-08 V_low
+ 2.080100000e-08 V_low
+ 2.090000000e-08 V_low
+ 2.090100000e-08 V_hig
+ 2.100000000e-08 V_hig
+ 2.100100000e-08 V_hig
+ 2.110000000e-08 V_hig
+ 2.110100000e-08 V_hig
+ 2.120000000e-08 V_hig
+ 2.120100000e-08 V_hig
+ 2.130000000e-08 V_hig
+ 2.130100000e-08 V_hig
+ 2.140000000e-08 V_hig
+ 2.140100000e-08 V_hig
+ 2.150000000e-08 V_hig
+ 2.150100000e-08 V_hig
+ 2.160000000e-08 V_hig
+ 2.160100000e-08 V_hig
+ 2.170000000e-08 V_hig
+ 2.170100000e-08 V_hig
+ 2.180000000e-08 V_hig
+ 2.180100000e-08 V_hig
+ 2.190000000e-08 V_hig
+ 2.190100000e-08 V_low
+ 2.200000000e-08 V_low
+ 2.200100000e-08 V_low
+ 2.210000000e-08 V_low
+ 2.210100000e-08 V_low
+ 2.220000000e-08 V_low
+ 2.220100000e-08 V_low
+ 2.230000000e-08 V_low
+ 2.230100000e-08 V_low
+ 2.240000000e-08 V_low
+ 2.240100000e-08 V_low
+ 2.250000000e-08 V_low
+ 2.250100000e-08 V_low
+ 2.260000000e-08 V_low
+ 2.260100000e-08 V_low
+ 2.270000000e-08 V_low
+ 2.270100000e-08 V_low
+ 2.280000000e-08 V_low
+ 2.280100000e-08 V_low
+ 2.290000000e-08 V_low
+ 2.290100000e-08 V_low
+ 2.300000000e-08 V_low
+ 2.300100000e-08 V_low
+ 2.310000000e-08 V_low
+ 2.310100000e-08 V_low
+ 2.320000000e-08 V_low
+ 2.320100000e-08 V_low
+ 2.330000000e-08 V_low
+ 2.330100000e-08 V_low
+ 2.340000000e-08 V_low
+ 2.340100000e-08 V_low
+ 2.350000000e-08 V_low
+ 2.350100000e-08 V_low
+ 2.360000000e-08 V_low
+ 2.360100000e-08 V_low
+ 2.370000000e-08 V_low
+ 2.370100000e-08 V_low
+ 2.380000000e-08 V_low
+ 2.380100000e-08 V_low
+ 2.390000000e-08 V_low
+ 2.390100000e-08 V_hig
+ 2.400000000e-08 V_hig
+ 2.400100000e-08 V_hig
+ 2.410000000e-08 V_hig
+ 2.410100000e-08 V_hig
+ 2.420000000e-08 V_hig
+ 2.420100000e-08 V_hig
+ 2.430000000e-08 V_hig
+ 2.430100000e-08 V_hig
+ 2.440000000e-08 V_hig
+ 2.440100000e-08 V_hig
+ 2.450000000e-08 V_hig
+ 2.450100000e-08 V_hig
+ 2.460000000e-08 V_hig
+ 2.460100000e-08 V_hig
+ 2.470000000e-08 V_hig
+ 2.470100000e-08 V_hig
+ 2.480000000e-08 V_hig
+ 2.480100000e-08 V_hig
+ 2.490000000e-08 V_hig
+ 2.490100000e-08 V_hig
+ 2.500000000e-08 V_hig
+ 2.500100000e-08 V_hig
+ 2.510000000e-08 V_hig
+ 2.510100000e-08 V_hig
+ 2.520000000e-08 V_hig
+ 2.520100000e-08 V_hig
+ 2.530000000e-08 V_hig
+ 2.530100000e-08 V_hig
+ 2.540000000e-08 V_hig
+ 2.540100000e-08 V_hig
+ 2.550000000e-08 V_hig
+ 2.550100000e-08 V_hig
+ 2.560000000e-08 V_hig
+ 2.560100000e-08 V_hig
+ 2.570000000e-08 V_hig
+ 2.570100000e-08 V_hig
+ 2.580000000e-08 V_hig
+ 2.580100000e-08 V_hig
+ 2.590000000e-08 V_hig
+ 2.590100000e-08 V_hig
+ 2.600000000e-08 V_hig
+ 2.600100000e-08 V_hig
+ 2.610000000e-08 V_hig
+ 2.610100000e-08 V_hig
+ 2.620000000e-08 V_hig
+ 2.620100000e-08 V_hig
+ 2.630000000e-08 V_hig
+ 2.630100000e-08 V_hig
+ 2.640000000e-08 V_hig
+ 2.640100000e-08 V_hig
+ 2.650000000e-08 V_hig
+ 2.650100000e-08 V_hig
+ 2.660000000e-08 V_hig
+ 2.660100000e-08 V_hig
+ 2.670000000e-08 V_hig
+ 2.670100000e-08 V_hig
+ 2.680000000e-08 V_hig
+ 2.680100000e-08 V_hig
+ 2.690000000e-08 V_hig
+ 2.690100000e-08 V_low
+ 2.700000000e-08 V_low
+ 2.700100000e-08 V_low
+ 2.710000000e-08 V_low
+ 2.710100000e-08 V_low
+ 2.720000000e-08 V_low
+ 2.720100000e-08 V_low
+ 2.730000000e-08 V_low
+ 2.730100000e-08 V_low
+ 2.740000000e-08 V_low
+ 2.740100000e-08 V_low
+ 2.750000000e-08 V_low
+ 2.750100000e-08 V_low
+ 2.760000000e-08 V_low
+ 2.760100000e-08 V_low
+ 2.770000000e-08 V_low
+ 2.770100000e-08 V_low
+ 2.780000000e-08 V_low
+ 2.780100000e-08 V_low
+ 2.790000000e-08 V_low
+ 2.790100000e-08 V_low
+ 2.800000000e-08 V_low
+ 2.800100000e-08 V_low
+ 2.810000000e-08 V_low
+ 2.810100000e-08 V_low
+ 2.820000000e-08 V_low
+ 2.820100000e-08 V_low
+ 2.830000000e-08 V_low
+ 2.830100000e-08 V_low
+ 2.840000000e-08 V_low
+ 2.840100000e-08 V_low
+ 2.850000000e-08 V_low
+ 2.850100000e-08 V_low
+ 2.860000000e-08 V_low
+ 2.860100000e-08 V_low
+ 2.870000000e-08 V_low
+ 2.870100000e-08 V_low
+ 2.880000000e-08 V_low
+ 2.880100000e-08 V_low
+ 2.890000000e-08 V_low
+ 2.890100000e-08 V_hig
+ 2.900000000e-08 V_hig
+ 2.900100000e-08 V_hig
+ 2.910000000e-08 V_hig
+ 2.910100000e-08 V_hig
+ 2.920000000e-08 V_hig
+ 2.920100000e-08 V_hig
+ 2.930000000e-08 V_hig
+ 2.930100000e-08 V_hig
+ 2.940000000e-08 V_hig
+ 2.940100000e-08 V_hig
+ 2.950000000e-08 V_hig
+ 2.950100000e-08 V_hig
+ 2.960000000e-08 V_hig
+ 2.960100000e-08 V_hig
+ 2.970000000e-08 V_hig
+ 2.970100000e-08 V_hig
+ 2.980000000e-08 V_hig
+ 2.980100000e-08 V_hig
+ 2.990000000e-08 V_hig
+ 2.990100000e-08 V_low
+ 3.000000000e-08 V_low
+ 3.000100000e-08 V_low
+ 3.010000000e-08 V_low
+ 3.010100000e-08 V_low
+ 3.020000000e-08 V_low
+ 3.020100000e-08 V_low
+ 3.030000000e-08 V_low
+ 3.030100000e-08 V_low
+ 3.040000000e-08 V_low
+ 3.040100000e-08 V_low
+ 3.050000000e-08 V_low
+ 3.050100000e-08 V_low
+ 3.060000000e-08 V_low
+ 3.060100000e-08 V_low
+ 3.070000000e-08 V_low
+ 3.070100000e-08 V_low
+ 3.080000000e-08 V_low
+ 3.080100000e-08 V_low
+ 3.090000000e-08 V_low
+ 3.090100000e-08 V_low
+ 3.100000000e-08 V_low
+ 3.100100000e-08 V_low
+ 3.110000000e-08 V_low
+ 3.110100000e-08 V_low
+ 3.120000000e-08 V_low
+ 3.120100000e-08 V_low
+ 3.130000000e-08 V_low
+ 3.130100000e-08 V_low
+ 3.140000000e-08 V_low
+ 3.140100000e-08 V_low
+ 3.150000000e-08 V_low
+ 3.150100000e-08 V_low
+ 3.160000000e-08 V_low
+ 3.160100000e-08 V_low
+ 3.170000000e-08 V_low
+ 3.170100000e-08 V_low
+ 3.180000000e-08 V_low
+ 3.180100000e-08 V_low
+ 3.190000000e-08 V_low
+ 3.190100000e-08 V_low
+ 3.200000000e-08 V_low
+ 3.200100000e-08 V_low
+ 3.210000000e-08 V_low
+ 3.210100000e-08 V_low
+ 3.220000000e-08 V_low
+ 3.220100000e-08 V_low
+ 3.230000000e-08 V_low
+ 3.230100000e-08 V_low
+ 3.240000000e-08 V_low
+ 3.240100000e-08 V_low
+ 3.250000000e-08 V_low
+ 3.250100000e-08 V_low
+ 3.260000000e-08 V_low
+ 3.260100000e-08 V_low
+ 3.270000000e-08 V_low
+ 3.270100000e-08 V_low
+ 3.280000000e-08 V_low
+ 3.280100000e-08 V_low
+ 3.290000000e-08 V_low
+ 3.290100000e-08 V_low
+ 3.300000000e-08 V_low
+ 3.300100000e-08 V_low
+ 3.310000000e-08 V_low
+ 3.310100000e-08 V_low
+ 3.320000000e-08 V_low
+ 3.320100000e-08 V_low
+ 3.330000000e-08 V_low
+ 3.330100000e-08 V_low
+ 3.340000000e-08 V_low
+ 3.340100000e-08 V_low
+ 3.350000000e-08 V_low
+ 3.350100000e-08 V_low
+ 3.360000000e-08 V_low
+ 3.360100000e-08 V_low
+ 3.370000000e-08 V_low
+ 3.370100000e-08 V_low
+ 3.380000000e-08 V_low
+ 3.380100000e-08 V_low
+ 3.390000000e-08 V_low
+ 3.390100000e-08 V_hig
+ 3.400000000e-08 V_hig
+ 3.400100000e-08 V_hig
+ 3.410000000e-08 V_hig
+ 3.410100000e-08 V_hig
+ 3.420000000e-08 V_hig
+ 3.420100000e-08 V_hig
+ 3.430000000e-08 V_hig
+ 3.430100000e-08 V_hig
+ 3.440000000e-08 V_hig
+ 3.440100000e-08 V_hig
+ 3.450000000e-08 V_hig
+ 3.450100000e-08 V_hig
+ 3.460000000e-08 V_hig
+ 3.460100000e-08 V_hig
+ 3.470000000e-08 V_hig
+ 3.470100000e-08 V_hig
+ 3.480000000e-08 V_hig
+ 3.480100000e-08 V_hig
+ 3.490000000e-08 V_hig
+ 3.490100000e-08 V_hig
+ 3.500000000e-08 V_hig
+ 3.500100000e-08 V_hig
+ 3.510000000e-08 V_hig
+ 3.510100000e-08 V_hig
+ 3.520000000e-08 V_hig
+ 3.520100000e-08 V_hig
+ 3.530000000e-08 V_hig
+ 3.530100000e-08 V_hig
+ 3.540000000e-08 V_hig
+ 3.540100000e-08 V_hig
+ 3.550000000e-08 V_hig
+ 3.550100000e-08 V_hig
+ 3.560000000e-08 V_hig
+ 3.560100000e-08 V_hig
+ 3.570000000e-08 V_hig
+ 3.570100000e-08 V_hig
+ 3.580000000e-08 V_hig
+ 3.580100000e-08 V_hig
+ 3.590000000e-08 V_hig
+ 3.590100000e-08 V_hig
+ 3.600000000e-08 V_hig
+ 3.600100000e-08 V_hig
+ 3.610000000e-08 V_hig
+ 3.610100000e-08 V_hig
+ 3.620000000e-08 V_hig
+ 3.620100000e-08 V_hig
+ 3.630000000e-08 V_hig
+ 3.630100000e-08 V_hig
+ 3.640000000e-08 V_hig
+ 3.640100000e-08 V_hig
+ 3.650000000e-08 V_hig
+ 3.650100000e-08 V_hig
+ 3.660000000e-08 V_hig
+ 3.660100000e-08 V_hig
+ 3.670000000e-08 V_hig
+ 3.670100000e-08 V_hig
+ 3.680000000e-08 V_hig
+ 3.680100000e-08 V_hig
+ 3.690000000e-08 V_hig
+ 3.690100000e-08 V_low
+ 3.700000000e-08 V_low
+ 3.700100000e-08 V_low
+ 3.710000000e-08 V_low
+ 3.710100000e-08 V_low
+ 3.720000000e-08 V_low
+ 3.720100000e-08 V_low
+ 3.730000000e-08 V_low
+ 3.730100000e-08 V_low
+ 3.740000000e-08 V_low
+ 3.740100000e-08 V_low
+ 3.750000000e-08 V_low
+ 3.750100000e-08 V_low
+ 3.760000000e-08 V_low
+ 3.760100000e-08 V_low
+ 3.770000000e-08 V_low
+ 3.770100000e-08 V_low
+ 3.780000000e-08 V_low
+ 3.780100000e-08 V_low
+ 3.790000000e-08 V_low
+ 3.790100000e-08 V_low
+ 3.800000000e-08 V_low
+ 3.800100000e-08 V_low
+ 3.810000000e-08 V_low
+ 3.810100000e-08 V_low
+ 3.820000000e-08 V_low
+ 3.820100000e-08 V_low
+ 3.830000000e-08 V_low
+ 3.830100000e-08 V_low
+ 3.840000000e-08 V_low
+ 3.840100000e-08 V_low
+ 3.850000000e-08 V_low
+ 3.850100000e-08 V_low
+ 3.860000000e-08 V_low
+ 3.860100000e-08 V_low
+ 3.870000000e-08 V_low
+ 3.870100000e-08 V_low
+ 3.880000000e-08 V_low
+ 3.880100000e-08 V_low
+ 3.890000000e-08 V_low
+ 3.890100000e-08 V_hig
+ 3.900000000e-08 V_hig
+ 3.900100000e-08 V_hig
+ 3.910000000e-08 V_hig
+ 3.910100000e-08 V_hig
+ 3.920000000e-08 V_hig
+ 3.920100000e-08 V_hig
+ 3.930000000e-08 V_hig
+ 3.930100000e-08 V_hig
+ 3.940000000e-08 V_hig
+ 3.940100000e-08 V_hig
+ 3.950000000e-08 V_hig
+ 3.950100000e-08 V_hig
+ 3.960000000e-08 V_hig
+ 3.960100000e-08 V_hig
+ 3.970000000e-08 V_hig
+ 3.970100000e-08 V_hig
+ 3.980000000e-08 V_hig
+ 3.980100000e-08 V_hig
+ 3.990000000e-08 V_hig
+ 3.990100000e-08 V_low
+ 4.000000000e-08 V_low
+ 4.000100000e-08 V_low
+ 4.010000000e-08 V_low
+ 4.010100000e-08 V_low
+ 4.020000000e-08 V_low
+ 4.020100000e-08 V_low
+ 4.030000000e-08 V_low
+ 4.030100000e-08 V_low
+ 4.040000000e-08 V_low
+ 4.040100000e-08 V_low
+ 4.050000000e-08 V_low
+ 4.050100000e-08 V_low
+ 4.060000000e-08 V_low
+ 4.060100000e-08 V_low
+ 4.070000000e-08 V_low
+ 4.070100000e-08 V_low
+ 4.080000000e-08 V_low
+ 4.080100000e-08 V_low
+ 4.090000000e-08 V_low
+ 4.090100000e-08 V_hig
+ 4.100000000e-08 V_hig
+ 4.100100000e-08 V_hig
+ 4.110000000e-08 V_hig
+ 4.110100000e-08 V_hig
+ 4.120000000e-08 V_hig
+ 4.120100000e-08 V_hig
+ 4.130000000e-08 V_hig
+ 4.130100000e-08 V_hig
+ 4.140000000e-08 V_hig
+ 4.140100000e-08 V_hig
+ 4.150000000e-08 V_hig
+ 4.150100000e-08 V_hig
+ 4.160000000e-08 V_hig
+ 4.160100000e-08 V_hig
+ 4.170000000e-08 V_hig
+ 4.170100000e-08 V_hig
+ 4.180000000e-08 V_hig
+ 4.180100000e-08 V_hig
+ 4.190000000e-08 V_hig
+ 4.190100000e-08 V_hig
+ 4.200000000e-08 V_hig
+ 4.200100000e-08 V_hig
+ 4.210000000e-08 V_hig
+ 4.210100000e-08 V_hig
+ 4.220000000e-08 V_hig
+ 4.220100000e-08 V_hig
+ 4.230000000e-08 V_hig
+ 4.230100000e-08 V_hig
+ 4.240000000e-08 V_hig
+ 4.240100000e-08 V_hig
+ 4.250000000e-08 V_hig
+ 4.250100000e-08 V_hig
+ 4.260000000e-08 V_hig
+ 4.260100000e-08 V_hig
+ 4.270000000e-08 V_hig
+ 4.270100000e-08 V_hig
+ 4.280000000e-08 V_hig
+ 4.280100000e-08 V_hig
+ 4.290000000e-08 V_hig
+ 4.290100000e-08 V_hig
+ 4.300000000e-08 V_hig
+ 4.300100000e-08 V_hig
+ 4.310000000e-08 V_hig
+ 4.310100000e-08 V_hig
+ 4.320000000e-08 V_hig
+ 4.320100000e-08 V_hig
+ 4.330000000e-08 V_hig
+ 4.330100000e-08 V_hig
+ 4.340000000e-08 V_hig
+ 4.340100000e-08 V_hig
+ 4.350000000e-08 V_hig
+ 4.350100000e-08 V_hig
+ 4.360000000e-08 V_hig
+ 4.360100000e-08 V_hig
+ 4.370000000e-08 V_hig
+ 4.370100000e-08 V_hig
+ 4.380000000e-08 V_hig
+ 4.380100000e-08 V_hig
+ 4.390000000e-08 V_hig
+ 4.390100000e-08 V_hig
+ 4.400000000e-08 V_hig
+ 4.400100000e-08 V_hig
+ 4.410000000e-08 V_hig
+ 4.410100000e-08 V_hig
+ 4.420000000e-08 V_hig
+ 4.420100000e-08 V_hig
+ 4.430000000e-08 V_hig
+ 4.430100000e-08 V_hig
+ 4.440000000e-08 V_hig
+ 4.440100000e-08 V_hig
+ 4.450000000e-08 V_hig
+ 4.450100000e-08 V_hig
+ 4.460000000e-08 V_hig
+ 4.460100000e-08 V_hig
+ 4.470000000e-08 V_hig
+ 4.470100000e-08 V_hig
+ 4.480000000e-08 V_hig
+ 4.480100000e-08 V_hig
+ 4.490000000e-08 V_hig
+ 4.490100000e-08 V_low
+ 4.500000000e-08 V_low
+ 4.500100000e-08 V_low
+ 4.510000000e-08 V_low
+ 4.510100000e-08 V_low
+ 4.520000000e-08 V_low
+ 4.520100000e-08 V_low
+ 4.530000000e-08 V_low
+ 4.530100000e-08 V_low
+ 4.540000000e-08 V_low
+ 4.540100000e-08 V_low
+ 4.550000000e-08 V_low
+ 4.550100000e-08 V_low
+ 4.560000000e-08 V_low
+ 4.560100000e-08 V_low
+ 4.570000000e-08 V_low
+ 4.570100000e-08 V_low
+ 4.580000000e-08 V_low
+ 4.580100000e-08 V_low
+ 4.590000000e-08 V_low
+ 4.590100000e-08 V_hig
+ 4.600000000e-08 V_hig
+ 4.600100000e-08 V_hig
+ 4.610000000e-08 V_hig
+ 4.610100000e-08 V_hig
+ 4.620000000e-08 V_hig
+ 4.620100000e-08 V_hig
+ 4.630000000e-08 V_hig
+ 4.630100000e-08 V_hig
+ 4.640000000e-08 V_hig
+ 4.640100000e-08 V_hig
+ 4.650000000e-08 V_hig
+ 4.650100000e-08 V_hig
+ 4.660000000e-08 V_hig
+ 4.660100000e-08 V_hig
+ 4.670000000e-08 V_hig
+ 4.670100000e-08 V_hig
+ 4.680000000e-08 V_hig
+ 4.680100000e-08 V_hig
+ 4.690000000e-08 V_hig
+ 4.690100000e-08 V_hig
+ 4.700000000e-08 V_hig
+ 4.700100000e-08 V_hig
+ 4.710000000e-08 V_hig
+ 4.710100000e-08 V_hig
+ 4.720000000e-08 V_hig
+ 4.720100000e-08 V_hig
+ 4.730000000e-08 V_hig
+ 4.730100000e-08 V_hig
+ 4.740000000e-08 V_hig
+ 4.740100000e-08 V_hig
+ 4.750000000e-08 V_hig
+ 4.750100000e-08 V_hig
+ 4.760000000e-08 V_hig
+ 4.760100000e-08 V_hig
+ 4.770000000e-08 V_hig
+ 4.770100000e-08 V_hig
+ 4.780000000e-08 V_hig
+ 4.780100000e-08 V_hig
+ 4.790000000e-08 V_hig
+ 4.790100000e-08 V_low
+ 4.800000000e-08 V_low
+ 4.800100000e-08 V_low
+ 4.810000000e-08 V_low
+ 4.810100000e-08 V_low
+ 4.820000000e-08 V_low
+ 4.820100000e-08 V_low
+ 4.830000000e-08 V_low
+ 4.830100000e-08 V_low
+ 4.840000000e-08 V_low
+ 4.840100000e-08 V_low
+ 4.850000000e-08 V_low
+ 4.850100000e-08 V_low
+ 4.860000000e-08 V_low
+ 4.860100000e-08 V_low
+ 4.870000000e-08 V_low
+ 4.870100000e-08 V_low
+ 4.880000000e-08 V_low
+ 4.880100000e-08 V_low
+ 4.890000000e-08 V_low
+ 4.890100000e-08 V_hig
+ 4.900000000e-08 V_hig
+ 4.900100000e-08 V_hig
+ 4.910000000e-08 V_hig
+ 4.910100000e-08 V_hig
+ 4.920000000e-08 V_hig
+ 4.920100000e-08 V_hig
+ 4.930000000e-08 V_hig
+ 4.930100000e-08 V_hig
+ 4.940000000e-08 V_hig
+ 4.940100000e-08 V_hig
+ 4.950000000e-08 V_hig
+ 4.950100000e-08 V_hig
+ 4.960000000e-08 V_hig
+ 4.960100000e-08 V_hig
+ 4.970000000e-08 V_hig
+ 4.970100000e-08 V_hig
+ 4.980000000e-08 V_hig
+ 4.980100000e-08 V_hig
+ 4.990000000e-08 V_hig
+ 4.990100000e-08 V_hig
+ 5.000000000e-08 V_hig
+ 5.000100000e-08 V_hig
+ 5.010000000e-08 V_hig
+ 5.010100000e-08 V_hig
+ 5.020000000e-08 V_hig
+ 5.020100000e-08 V_hig
+ 5.030000000e-08 V_hig
+ 5.030100000e-08 V_hig
+ 5.040000000e-08 V_hig
+ 5.040100000e-08 V_hig
+ 5.050000000e-08 V_hig
+ 5.050100000e-08 V_hig
+ 5.060000000e-08 V_hig
+ 5.060100000e-08 V_hig
+ 5.070000000e-08 V_hig
+ 5.070100000e-08 V_hig
+ 5.080000000e-08 V_hig
+ 5.080100000e-08 V_hig
+ 5.090000000e-08 V_hig
+ 5.090100000e-08 V_hig
+ 5.100000000e-08 V_hig
+ 5.100100000e-08 V_hig
+ 5.110000000e-08 V_hig
+ 5.110100000e-08 V_hig
+ 5.120000000e-08 V_hig
+ 5.120100000e-08 V_hig
+ 5.130000000e-08 V_hig
+ 5.130100000e-08 V_hig
+ 5.140000000e-08 V_hig
+ 5.140100000e-08 V_hig
+ 5.150000000e-08 V_hig
+ 5.150100000e-08 V_hig
+ 5.160000000e-08 V_hig
+ 5.160100000e-08 V_hig
+ 5.170000000e-08 V_hig
+ 5.170100000e-08 V_hig
+ 5.180000000e-08 V_hig
+ 5.180100000e-08 V_hig
+ 5.190000000e-08 V_hig
+ 5.190100000e-08 V_low
+ 5.200000000e-08 V_low
+ 5.200100000e-08 V_low
+ 5.210000000e-08 V_low
+ 5.210100000e-08 V_low
+ 5.220000000e-08 V_low
+ 5.220100000e-08 V_low
+ 5.230000000e-08 V_low
+ 5.230100000e-08 V_low
+ 5.240000000e-08 V_low
+ 5.240100000e-08 V_low
+ 5.250000000e-08 V_low
+ 5.250100000e-08 V_low
+ 5.260000000e-08 V_low
+ 5.260100000e-08 V_low
+ 5.270000000e-08 V_low
+ 5.270100000e-08 V_low
+ 5.280000000e-08 V_low
+ 5.280100000e-08 V_low
+ 5.290000000e-08 V_low
+ 5.290100000e-08 V_low
+ 5.300000000e-08 V_low
+ 5.300100000e-08 V_low
+ 5.310000000e-08 V_low
+ 5.310100000e-08 V_low
+ 5.320000000e-08 V_low
+ 5.320100000e-08 V_low
+ 5.330000000e-08 V_low
+ 5.330100000e-08 V_low
+ 5.340000000e-08 V_low
+ 5.340100000e-08 V_low
+ 5.350000000e-08 V_low
+ 5.350100000e-08 V_low
+ 5.360000000e-08 V_low
+ 5.360100000e-08 V_low
+ 5.370000000e-08 V_low
+ 5.370100000e-08 V_low
+ 5.380000000e-08 V_low
+ 5.380100000e-08 V_low
+ 5.390000000e-08 V_low
+ 5.390100000e-08 V_hig
+ 5.400000000e-08 V_hig
+ 5.400100000e-08 V_hig
+ 5.410000000e-08 V_hig
+ 5.410100000e-08 V_hig
+ 5.420000000e-08 V_hig
+ 5.420100000e-08 V_hig
+ 5.430000000e-08 V_hig
+ 5.430100000e-08 V_hig
+ 5.440000000e-08 V_hig
+ 5.440100000e-08 V_hig
+ 5.450000000e-08 V_hig
+ 5.450100000e-08 V_hig
+ 5.460000000e-08 V_hig
+ 5.460100000e-08 V_hig
+ 5.470000000e-08 V_hig
+ 5.470100000e-08 V_hig
+ 5.480000000e-08 V_hig
+ 5.480100000e-08 V_hig
+ 5.490000000e-08 V_hig
+ 5.490100000e-08 V_low
+ 5.500000000e-08 V_low
+ 5.500100000e-08 V_low
+ 5.510000000e-08 V_low
+ 5.510100000e-08 V_low
+ 5.520000000e-08 V_low
+ 5.520100000e-08 V_low
+ 5.530000000e-08 V_low
+ 5.530100000e-08 V_low
+ 5.540000000e-08 V_low
+ 5.540100000e-08 V_low
+ 5.550000000e-08 V_low
+ 5.550100000e-08 V_low
+ 5.560000000e-08 V_low
+ 5.560100000e-08 V_low
+ 5.570000000e-08 V_low
+ 5.570100000e-08 V_low
+ 5.580000000e-08 V_low
+ 5.580100000e-08 V_low
+ 5.590000000e-08 V_low
+ 5.590100000e-08 V_hig
+ 5.600000000e-08 V_hig
+ 5.600100000e-08 V_hig
+ 5.610000000e-08 V_hig
+ 5.610100000e-08 V_hig
+ 5.620000000e-08 V_hig
+ 5.620100000e-08 V_hig
+ 5.630000000e-08 V_hig
+ 5.630100000e-08 V_hig
+ 5.640000000e-08 V_hig
+ 5.640100000e-08 V_hig
+ 5.650000000e-08 V_hig
+ 5.650100000e-08 V_hig
+ 5.660000000e-08 V_hig
+ 5.660100000e-08 V_hig
+ 5.670000000e-08 V_hig
+ 5.670100000e-08 V_hig
+ 5.680000000e-08 V_hig
+ 5.680100000e-08 V_hig
+ 5.690000000e-08 V_hig
+ 5.690100000e-08 V_low
+ 5.700000000e-08 V_low
+ 5.700100000e-08 V_low
+ 5.710000000e-08 V_low
+ 5.710100000e-08 V_low
+ 5.720000000e-08 V_low
+ 5.720100000e-08 V_low
+ 5.730000000e-08 V_low
+ 5.730100000e-08 V_low
+ 5.740000000e-08 V_low
+ 5.740100000e-08 V_low
+ 5.750000000e-08 V_low
+ 5.750100000e-08 V_low
+ 5.760000000e-08 V_low
+ 5.760100000e-08 V_low
+ 5.770000000e-08 V_low
+ 5.770100000e-08 V_low
+ 5.780000000e-08 V_low
+ 5.780100000e-08 V_low
+ 5.790000000e-08 V_low
+ 5.790100000e-08 V_hig
+ 5.800000000e-08 V_hig
+ 5.800100000e-08 V_hig
+ 5.810000000e-08 V_hig
+ 5.810100000e-08 V_hig
+ 5.820000000e-08 V_hig
+ 5.820100000e-08 V_hig
+ 5.830000000e-08 V_hig
+ 5.830100000e-08 V_hig
+ 5.840000000e-08 V_hig
+ 5.840100000e-08 V_hig
+ 5.850000000e-08 V_hig
+ 5.850100000e-08 V_hig
+ 5.860000000e-08 V_hig
+ 5.860100000e-08 V_hig
+ 5.870000000e-08 V_hig
+ 5.870100000e-08 V_hig
+ 5.880000000e-08 V_hig
+ 5.880100000e-08 V_hig
+ 5.890000000e-08 V_hig
+ 5.890100000e-08 V_low
+ 5.900000000e-08 V_low
+ 5.900100000e-08 V_low
+ 5.910000000e-08 V_low
+ 5.910100000e-08 V_low
+ 5.920000000e-08 V_low
+ 5.920100000e-08 V_low
+ 5.930000000e-08 V_low
+ 5.930100000e-08 V_low
+ 5.940000000e-08 V_low
+ 5.940100000e-08 V_low
+ 5.950000000e-08 V_low
+ 5.950100000e-08 V_low
+ 5.960000000e-08 V_low
+ 5.960100000e-08 V_low
+ 5.970000000e-08 V_low
+ 5.970100000e-08 V_low
+ 5.980000000e-08 V_low
+ 5.980100000e-08 V_low
+ 5.990000000e-08 V_low
+ 5.990100000e-08 V_hig
+ 6.000000000e-08 V_hig
+ 6.000100000e-08 V_hig
+ 6.010000000e-08 V_hig
+ 6.010100000e-08 V_hig
+ 6.020000000e-08 V_hig
+ 6.020100000e-08 V_hig
+ 6.030000000e-08 V_hig
+ 6.030100000e-08 V_hig
+ 6.040000000e-08 V_hig
+ 6.040100000e-08 V_hig
+ 6.050000000e-08 V_hig
+ 6.050100000e-08 V_hig
+ 6.060000000e-08 V_hig
+ 6.060100000e-08 V_hig
+ 6.070000000e-08 V_hig
+ 6.070100000e-08 V_hig
+ 6.080000000e-08 V_hig
+ 6.080100000e-08 V_hig
+ 6.090000000e-08 V_hig
+ 6.090100000e-08 V_hig
+ 6.100000000e-08 V_hig
+ 6.100100000e-08 V_hig
+ 6.110000000e-08 V_hig
+ 6.110100000e-08 V_hig
+ 6.120000000e-08 V_hig
+ 6.120100000e-08 V_hig
+ 6.130000000e-08 V_hig
+ 6.130100000e-08 V_hig
+ 6.140000000e-08 V_hig
+ 6.140100000e-08 V_hig
+ 6.150000000e-08 V_hig
+ 6.150100000e-08 V_hig
+ 6.160000000e-08 V_hig
+ 6.160100000e-08 V_hig
+ 6.170000000e-08 V_hig
+ 6.170100000e-08 V_hig
+ 6.180000000e-08 V_hig
+ 6.180100000e-08 V_hig
+ 6.190000000e-08 V_hig
+ 6.190100000e-08 V_hig
+ 6.200000000e-08 V_hig
+ 6.200100000e-08 V_hig
+ 6.210000000e-08 V_hig
+ 6.210100000e-08 V_hig
+ 6.220000000e-08 V_hig
+ 6.220100000e-08 V_hig
+ 6.230000000e-08 V_hig
+ 6.230100000e-08 V_hig
+ 6.240000000e-08 V_hig
+ 6.240100000e-08 V_hig
+ 6.250000000e-08 V_hig
+ 6.250100000e-08 V_hig
+ 6.260000000e-08 V_hig
+ 6.260100000e-08 V_hig
+ 6.270000000e-08 V_hig
+ 6.270100000e-08 V_hig
+ 6.280000000e-08 V_hig
+ 6.280100000e-08 V_hig
+ 6.290000000e-08 V_hig
+ 6.290100000e-08 V_hig
+ 6.300000000e-08 V_hig
+ 6.300100000e-08 V_hig
+ 6.310000000e-08 V_hig
+ 6.310100000e-08 V_hig
+ 6.320000000e-08 V_hig
+ 6.320100000e-08 V_hig
+ 6.330000000e-08 V_hig
+ 6.330100000e-08 V_hig
+ 6.340000000e-08 V_hig
+ 6.340100000e-08 V_hig
+ 6.350000000e-08 V_hig
+ 6.350100000e-08 V_hig
+ 6.360000000e-08 V_hig
+ 6.360100000e-08 V_hig
+ 6.370000000e-08 V_hig
+ 6.370100000e-08 V_hig
+ 6.380000000e-08 V_hig
+ 6.380100000e-08 V_hig
+ 6.390000000e-08 V_hig
+ 6.390100000e-08 V_hig
+ 6.400000000e-08 V_hig
+ 6.400100000e-08 V_hig
+ 6.410000000e-08 V_hig
+ 6.410100000e-08 V_hig
+ 6.420000000e-08 V_hig
+ 6.420100000e-08 V_hig
+ 6.430000000e-08 V_hig
+ 6.430100000e-08 V_hig
+ 6.440000000e-08 V_hig
+ 6.440100000e-08 V_hig
+ 6.450000000e-08 V_hig
+ 6.450100000e-08 V_hig
+ 6.460000000e-08 V_hig
+ 6.460100000e-08 V_hig
+ 6.470000000e-08 V_hig
+ 6.470100000e-08 V_hig
+ 6.480000000e-08 V_hig
+ 6.480100000e-08 V_hig
+ 6.490000000e-08 V_hig
+ 6.490100000e-08 V_hig
+ 6.500000000e-08 V_hig
+ 6.500100000e-08 V_hig
+ 6.510000000e-08 V_hig
+ 6.510100000e-08 V_hig
+ 6.520000000e-08 V_hig
+ 6.520100000e-08 V_hig
+ 6.530000000e-08 V_hig
+ 6.530100000e-08 V_hig
+ 6.540000000e-08 V_hig
+ 6.540100000e-08 V_hig
+ 6.550000000e-08 V_hig
+ 6.550100000e-08 V_hig
+ 6.560000000e-08 V_hig
+ 6.560100000e-08 V_hig
+ 6.570000000e-08 V_hig
+ 6.570100000e-08 V_hig
+ 6.580000000e-08 V_hig
+ 6.580100000e-08 V_hig
+ 6.590000000e-08 V_hig
+ 6.590100000e-08 V_hig
+ 6.600000000e-08 V_hig
+ 6.600100000e-08 V_hig
+ 6.610000000e-08 V_hig
+ 6.610100000e-08 V_hig
+ 6.620000000e-08 V_hig
+ 6.620100000e-08 V_hig
+ 6.630000000e-08 V_hig
+ 6.630100000e-08 V_hig
+ 6.640000000e-08 V_hig
+ 6.640100000e-08 V_hig
+ 6.650000000e-08 V_hig
+ 6.650100000e-08 V_hig
+ 6.660000000e-08 V_hig
+ 6.660100000e-08 V_hig
+ 6.670000000e-08 V_hig
+ 6.670100000e-08 V_hig
+ 6.680000000e-08 V_hig
+ 6.680100000e-08 V_hig
+ 6.690000000e-08 V_hig
+ 6.690100000e-08 V_low
+ 6.700000000e-08 V_low
+ 6.700100000e-08 V_low
+ 6.710000000e-08 V_low
+ 6.710100000e-08 V_low
+ 6.720000000e-08 V_low
+ 6.720100000e-08 V_low
+ 6.730000000e-08 V_low
+ 6.730100000e-08 V_low
+ 6.740000000e-08 V_low
+ 6.740100000e-08 V_low
+ 6.750000000e-08 V_low
+ 6.750100000e-08 V_low
+ 6.760000000e-08 V_low
+ 6.760100000e-08 V_low
+ 6.770000000e-08 V_low
+ 6.770100000e-08 V_low
+ 6.780000000e-08 V_low
+ 6.780100000e-08 V_low
+ 6.790000000e-08 V_low
+ 6.790100000e-08 V_low
+ 6.800000000e-08 V_low
+ 6.800100000e-08 V_low
+ 6.810000000e-08 V_low
+ 6.810100000e-08 V_low
+ 6.820000000e-08 V_low
+ 6.820100000e-08 V_low
+ 6.830000000e-08 V_low
+ 6.830100000e-08 V_low
+ 6.840000000e-08 V_low
+ 6.840100000e-08 V_low
+ 6.850000000e-08 V_low
+ 6.850100000e-08 V_low
+ 6.860000000e-08 V_low
+ 6.860100000e-08 V_low
+ 6.870000000e-08 V_low
+ 6.870100000e-08 V_low
+ 6.880000000e-08 V_low
+ 6.880100000e-08 V_low
+ 6.890000000e-08 V_low
+ 6.890100000e-08 V_hig
+ 6.900000000e-08 V_hig
+ 6.900100000e-08 V_hig
+ 6.910000000e-08 V_hig
+ 6.910100000e-08 V_hig
+ 6.920000000e-08 V_hig
+ 6.920100000e-08 V_hig
+ 6.930000000e-08 V_hig
+ 6.930100000e-08 V_hig
+ 6.940000000e-08 V_hig
+ 6.940100000e-08 V_hig
+ 6.950000000e-08 V_hig
+ 6.950100000e-08 V_hig
+ 6.960000000e-08 V_hig
+ 6.960100000e-08 V_hig
+ 6.970000000e-08 V_hig
+ 6.970100000e-08 V_hig
+ 6.980000000e-08 V_hig
+ 6.980100000e-08 V_hig
+ 6.990000000e-08 V_hig
+ 6.990100000e-08 V_hig
+ 7.000000000e-08 V_hig
+ 7.000100000e-08 V_hig
+ 7.010000000e-08 V_hig
+ 7.010100000e-08 V_hig
+ 7.020000000e-08 V_hig
+ 7.020100000e-08 V_hig
+ 7.030000000e-08 V_hig
+ 7.030100000e-08 V_hig
+ 7.040000000e-08 V_hig
+ 7.040100000e-08 V_hig
+ 7.050000000e-08 V_hig
+ 7.050100000e-08 V_hig
+ 7.060000000e-08 V_hig
+ 7.060100000e-08 V_hig
+ 7.070000000e-08 V_hig
+ 7.070100000e-08 V_hig
+ 7.080000000e-08 V_hig
+ 7.080100000e-08 V_hig
+ 7.090000000e-08 V_hig
+ 7.090100000e-08 V_hig
+ 7.100000000e-08 V_hig
+ 7.100100000e-08 V_hig
+ 7.110000000e-08 V_hig
+ 7.110100000e-08 V_hig
+ 7.120000000e-08 V_hig
+ 7.120100000e-08 V_hig
+ 7.130000000e-08 V_hig
+ 7.130100000e-08 V_hig
+ 7.140000000e-08 V_hig
+ 7.140100000e-08 V_hig
+ 7.150000000e-08 V_hig
+ 7.150100000e-08 V_hig
+ 7.160000000e-08 V_hig
+ 7.160100000e-08 V_hig
+ 7.170000000e-08 V_hig
+ 7.170100000e-08 V_hig
+ 7.180000000e-08 V_hig
+ 7.180100000e-08 V_hig
+ 7.190000000e-08 V_hig
+ 7.190100000e-08 V_hig
+ 7.200000000e-08 V_hig
+ 7.200100000e-08 V_hig
+ 7.210000000e-08 V_hig
+ 7.210100000e-08 V_hig
+ 7.220000000e-08 V_hig
+ 7.220100000e-08 V_hig
+ 7.230000000e-08 V_hig
+ 7.230100000e-08 V_hig
+ 7.240000000e-08 V_hig
+ 7.240100000e-08 V_hig
+ 7.250000000e-08 V_hig
+ 7.250100000e-08 V_hig
+ 7.260000000e-08 V_hig
+ 7.260100000e-08 V_hig
+ 7.270000000e-08 V_hig
+ 7.270100000e-08 V_hig
+ 7.280000000e-08 V_hig
+ 7.280100000e-08 V_hig
+ 7.290000000e-08 V_hig
+ 7.290100000e-08 V_hig
+ 7.300000000e-08 V_hig
+ 7.300100000e-08 V_hig
+ 7.310000000e-08 V_hig
+ 7.310100000e-08 V_hig
+ 7.320000000e-08 V_hig
+ 7.320100000e-08 V_hig
+ 7.330000000e-08 V_hig
+ 7.330100000e-08 V_hig
+ 7.340000000e-08 V_hig
+ 7.340100000e-08 V_hig
+ 7.350000000e-08 V_hig
+ 7.350100000e-08 V_hig
+ 7.360000000e-08 V_hig
+ 7.360100000e-08 V_hig
+ 7.370000000e-08 V_hig
+ 7.370100000e-08 V_hig
+ 7.380000000e-08 V_hig
+ 7.380100000e-08 V_hig
+ 7.390000000e-08 V_hig
+ 7.390100000e-08 V_hig
+ 7.400000000e-08 V_hig
+ 7.400100000e-08 V_hig
+ 7.410000000e-08 V_hig
+ 7.410100000e-08 V_hig
+ 7.420000000e-08 V_hig
+ 7.420100000e-08 V_hig
+ 7.430000000e-08 V_hig
+ 7.430100000e-08 V_hig
+ 7.440000000e-08 V_hig
+ 7.440100000e-08 V_hig
+ 7.450000000e-08 V_hig
+ 7.450100000e-08 V_hig
+ 7.460000000e-08 V_hig
+ 7.460100000e-08 V_hig
+ 7.470000000e-08 V_hig
+ 7.470100000e-08 V_hig
+ 7.480000000e-08 V_hig
+ 7.480100000e-08 V_hig
+ 7.490000000e-08 V_hig
+ 7.490100000e-08 V_low
+ 7.500000000e-08 V_low
+ 7.500100000e-08 V_low
+ 7.510000000e-08 V_low
+ 7.510100000e-08 V_low
+ 7.520000000e-08 V_low
+ 7.520100000e-08 V_low
+ 7.530000000e-08 V_low
+ 7.530100000e-08 V_low
+ 7.540000000e-08 V_low
+ 7.540100000e-08 V_low
+ 7.550000000e-08 V_low
+ 7.550100000e-08 V_low
+ 7.560000000e-08 V_low
+ 7.560100000e-08 V_low
+ 7.570000000e-08 V_low
+ 7.570100000e-08 V_low
+ 7.580000000e-08 V_low
+ 7.580100000e-08 V_low
+ 7.590000000e-08 V_low
+ 7.590100000e-08 V_low
+ 7.600000000e-08 V_low
+ 7.600100000e-08 V_low
+ 7.610000000e-08 V_low
+ 7.610100000e-08 V_low
+ 7.620000000e-08 V_low
+ 7.620100000e-08 V_low
+ 7.630000000e-08 V_low
+ 7.630100000e-08 V_low
+ 7.640000000e-08 V_low
+ 7.640100000e-08 V_low
+ 7.650000000e-08 V_low
+ 7.650100000e-08 V_low
+ 7.660000000e-08 V_low
+ 7.660100000e-08 V_low
+ 7.670000000e-08 V_low
+ 7.670100000e-08 V_low
+ 7.680000000e-08 V_low
+ 7.680100000e-08 V_low
+ 7.690000000e-08 V_low
+ 7.690100000e-08 V_hig
+ 7.700000000e-08 V_hig
+ 7.700100000e-08 V_hig
+ 7.710000000e-08 V_hig
+ 7.710100000e-08 V_hig
+ 7.720000000e-08 V_hig
+ 7.720100000e-08 V_hig
+ 7.730000000e-08 V_hig
+ 7.730100000e-08 V_hig
+ 7.740000000e-08 V_hig
+ 7.740100000e-08 V_hig
+ 7.750000000e-08 V_hig
+ 7.750100000e-08 V_hig
+ 7.760000000e-08 V_hig
+ 7.760100000e-08 V_hig
+ 7.770000000e-08 V_hig
+ 7.770100000e-08 V_hig
+ 7.780000000e-08 V_hig
+ 7.780100000e-08 V_hig
+ 7.790000000e-08 V_hig
+ 7.790100000e-08 V_hig
+ 7.800000000e-08 V_hig
+ 7.800100000e-08 V_hig
+ 7.810000000e-08 V_hig
+ 7.810100000e-08 V_hig
+ 7.820000000e-08 V_hig
+ 7.820100000e-08 V_hig
+ 7.830000000e-08 V_hig
+ 7.830100000e-08 V_hig
+ 7.840000000e-08 V_hig
+ 7.840100000e-08 V_hig
+ 7.850000000e-08 V_hig
+ 7.850100000e-08 V_hig
+ 7.860000000e-08 V_hig
+ 7.860100000e-08 V_hig
+ 7.870000000e-08 V_hig
+ 7.870100000e-08 V_hig
+ 7.880000000e-08 V_hig
+ 7.880100000e-08 V_hig
+ 7.890000000e-08 V_hig
+ 7.890100000e-08 V_low
+ 7.900000000e-08 V_low
+ 7.900100000e-08 V_low
+ 7.910000000e-08 V_low
+ 7.910100000e-08 V_low
+ 7.920000000e-08 V_low
+ 7.920100000e-08 V_low
+ 7.930000000e-08 V_low
+ 7.930100000e-08 V_low
+ 7.940000000e-08 V_low
+ 7.940100000e-08 V_low
+ 7.950000000e-08 V_low
+ 7.950100000e-08 V_low
+ 7.960000000e-08 V_low
+ 7.960100000e-08 V_low
+ 7.970000000e-08 V_low
+ 7.970100000e-08 V_low
+ 7.980000000e-08 V_low
+ 7.980100000e-08 V_low
+ 7.990000000e-08 V_low
+ 7.990100000e-08 V_low
+ 8.000000000e-08 V_low
+ 8.000100000e-08 V_low
+ 8.010000000e-08 V_low
+ 8.010100000e-08 V_low
+ 8.020000000e-08 V_low
+ 8.020100000e-08 V_low
+ 8.030000000e-08 V_low
+ 8.030100000e-08 V_low
+ 8.040000000e-08 V_low
+ 8.040100000e-08 V_low
+ 8.050000000e-08 V_low
+ 8.050100000e-08 V_low
+ 8.060000000e-08 V_low
+ 8.060100000e-08 V_low
+ 8.070000000e-08 V_low
+ 8.070100000e-08 V_low
+ 8.080000000e-08 V_low
+ 8.080100000e-08 V_low
+ 8.090000000e-08 V_low
+ 8.090100000e-08 V_hig
+ 8.100000000e-08 V_hig
+ 8.100100000e-08 V_hig
+ 8.110000000e-08 V_hig
+ 8.110100000e-08 V_hig
+ 8.120000000e-08 V_hig
+ 8.120100000e-08 V_hig
+ 8.130000000e-08 V_hig
+ 8.130100000e-08 V_hig
+ 8.140000000e-08 V_hig
+ 8.140100000e-08 V_hig
+ 8.150000000e-08 V_hig
+ 8.150100000e-08 V_hig
+ 8.160000000e-08 V_hig
+ 8.160100000e-08 V_hig
+ 8.170000000e-08 V_hig
+ 8.170100000e-08 V_hig
+ 8.180000000e-08 V_hig
+ 8.180100000e-08 V_hig
+ 8.190000000e-08 V_hig
+ 8.190100000e-08 V_hig
+ 8.200000000e-08 V_hig
+ 8.200100000e-08 V_hig
+ 8.210000000e-08 V_hig
+ 8.210100000e-08 V_hig
+ 8.220000000e-08 V_hig
+ 8.220100000e-08 V_hig
+ 8.230000000e-08 V_hig
+ 8.230100000e-08 V_hig
+ 8.240000000e-08 V_hig
+ 8.240100000e-08 V_hig
+ 8.250000000e-08 V_hig
+ 8.250100000e-08 V_hig
+ 8.260000000e-08 V_hig
+ 8.260100000e-08 V_hig
+ 8.270000000e-08 V_hig
+ 8.270100000e-08 V_hig
+ 8.280000000e-08 V_hig
+ 8.280100000e-08 V_hig
+ 8.290000000e-08 V_hig
+ 8.290100000e-08 V_hig
+ 8.300000000e-08 V_hig
+ 8.300100000e-08 V_hig
+ 8.310000000e-08 V_hig
+ 8.310100000e-08 V_hig
+ 8.320000000e-08 V_hig
+ 8.320100000e-08 V_hig
+ 8.330000000e-08 V_hig
+ 8.330100000e-08 V_hig
+ 8.340000000e-08 V_hig
+ 8.340100000e-08 V_hig
+ 8.350000000e-08 V_hig
+ 8.350100000e-08 V_hig
+ 8.360000000e-08 V_hig
+ 8.360100000e-08 V_hig
+ 8.370000000e-08 V_hig
+ 8.370100000e-08 V_hig
+ 8.380000000e-08 V_hig
+ 8.380100000e-08 V_hig
+ 8.390000000e-08 V_hig
+ 8.390100000e-08 V_low
+ 8.400000000e-08 V_low
+ 8.400100000e-08 V_low
+ 8.410000000e-08 V_low
+ 8.410100000e-08 V_low
+ 8.420000000e-08 V_low
+ 8.420100000e-08 V_low
+ 8.430000000e-08 V_low
+ 8.430100000e-08 V_low
+ 8.440000000e-08 V_low
+ 8.440100000e-08 V_low
+ 8.450000000e-08 V_low
+ 8.450100000e-08 V_low
+ 8.460000000e-08 V_low
+ 8.460100000e-08 V_low
+ 8.470000000e-08 V_low
+ 8.470100000e-08 V_low
+ 8.480000000e-08 V_low
+ 8.480100000e-08 V_low
+ 8.490000000e-08 V_low
+ 8.490100000e-08 V_hig
+ 8.500000000e-08 V_hig
+ 8.500100000e-08 V_hig
+ 8.510000000e-08 V_hig
+ 8.510100000e-08 V_hig
+ 8.520000000e-08 V_hig
+ 8.520100000e-08 V_hig
+ 8.530000000e-08 V_hig
+ 8.530100000e-08 V_hig
+ 8.540000000e-08 V_hig
+ 8.540100000e-08 V_hig
+ 8.550000000e-08 V_hig
+ 8.550100000e-08 V_hig
+ 8.560000000e-08 V_hig
+ 8.560100000e-08 V_hig
+ 8.570000000e-08 V_hig
+ 8.570100000e-08 V_hig
+ 8.580000000e-08 V_hig
+ 8.580100000e-08 V_hig
+ 8.590000000e-08 V_hig
+ 8.590100000e-08 V_low
+ 8.600000000e-08 V_low
+ 8.600100000e-08 V_low
+ 8.610000000e-08 V_low
+ 8.610100000e-08 V_low
+ 8.620000000e-08 V_low
+ 8.620100000e-08 V_low
+ 8.630000000e-08 V_low
+ 8.630100000e-08 V_low
+ 8.640000000e-08 V_low
+ 8.640100000e-08 V_low
+ 8.650000000e-08 V_low
+ 8.650100000e-08 V_low
+ 8.660000000e-08 V_low
+ 8.660100000e-08 V_low
+ 8.670000000e-08 V_low
+ 8.670100000e-08 V_low
+ 8.680000000e-08 V_low
+ 8.680100000e-08 V_low
+ 8.690000000e-08 V_low
+ 8.690100000e-08 V_low
+ 8.700000000e-08 V_low
+ 8.700100000e-08 V_low
+ 8.710000000e-08 V_low
+ 8.710100000e-08 V_low
+ 8.720000000e-08 V_low
+ 8.720100000e-08 V_low
+ 8.730000000e-08 V_low
+ 8.730100000e-08 V_low
+ 8.740000000e-08 V_low
+ 8.740100000e-08 V_low
+ 8.750000000e-08 V_low
+ 8.750100000e-08 V_low
+ 8.760000000e-08 V_low
+ 8.760100000e-08 V_low
+ 8.770000000e-08 V_low
+ 8.770100000e-08 V_low
+ 8.780000000e-08 V_low
+ 8.780100000e-08 V_low
+ 8.790000000e-08 V_low
+ 8.790100000e-08 V_hig
+ 8.800000000e-08 V_hig
+ 8.800100000e-08 V_hig
+ 8.810000000e-08 V_hig
+ 8.810100000e-08 V_hig
+ 8.820000000e-08 V_hig
+ 8.820100000e-08 V_hig
+ 8.830000000e-08 V_hig
+ 8.830100000e-08 V_hig
+ 8.840000000e-08 V_hig
+ 8.840100000e-08 V_hig
+ 8.850000000e-08 V_hig
+ 8.850100000e-08 V_hig
+ 8.860000000e-08 V_hig
+ 8.860100000e-08 V_hig
+ 8.870000000e-08 V_hig
+ 8.870100000e-08 V_hig
+ 8.880000000e-08 V_hig
+ 8.880100000e-08 V_hig
+ 8.890000000e-08 V_hig
+ 8.890100000e-08 V_low
+ 8.900000000e-08 V_low
+ 8.900100000e-08 V_low
+ 8.910000000e-08 V_low
+ 8.910100000e-08 V_low
+ 8.920000000e-08 V_low
+ 8.920100000e-08 V_low
+ 8.930000000e-08 V_low
+ 8.930100000e-08 V_low
+ 8.940000000e-08 V_low
+ 8.940100000e-08 V_low
+ 8.950000000e-08 V_low
+ 8.950100000e-08 V_low
+ 8.960000000e-08 V_low
+ 8.960100000e-08 V_low
+ 8.970000000e-08 V_low
+ 8.970100000e-08 V_low
+ 8.980000000e-08 V_low
+ 8.980100000e-08 V_low
+ 8.990000000e-08 V_low
+ 8.990100000e-08 V_low
+ 9.000000000e-08 V_low
+ 9.000100000e-08 V_low
+ 9.010000000e-08 V_low
+ 9.010100000e-08 V_low
+ 9.020000000e-08 V_low
+ 9.020100000e-08 V_low
+ 9.030000000e-08 V_low
+ 9.030100000e-08 V_low
+ 9.040000000e-08 V_low
+ 9.040100000e-08 V_low
+ 9.050000000e-08 V_low
+ 9.050100000e-08 V_low
+ 9.060000000e-08 V_low
+ 9.060100000e-08 V_low
+ 9.070000000e-08 V_low
+ 9.070100000e-08 V_low
+ 9.080000000e-08 V_low
+ 9.080100000e-08 V_low
+ 9.090000000e-08 V_low
+ 9.090100000e-08 V_low
+ 9.100000000e-08 V_low
+ 9.100100000e-08 V_low
+ 9.110000000e-08 V_low
+ 9.110100000e-08 V_low
+ 9.120000000e-08 V_low
+ 9.120100000e-08 V_low
+ 9.130000000e-08 V_low
+ 9.130100000e-08 V_low
+ 9.140000000e-08 V_low
+ 9.140100000e-08 V_low
+ 9.150000000e-08 V_low
+ 9.150100000e-08 V_low
+ 9.160000000e-08 V_low
+ 9.160100000e-08 V_low
+ 9.170000000e-08 V_low
+ 9.170100000e-08 V_low
+ 9.180000000e-08 V_low
+ 9.180100000e-08 V_low
+ 9.190000000e-08 V_low
+ 9.190100000e-08 V_hig
+ 9.200000000e-08 V_hig
+ 9.200100000e-08 V_hig
+ 9.210000000e-08 V_hig
+ 9.210100000e-08 V_hig
+ 9.220000000e-08 V_hig
+ 9.220100000e-08 V_hig
+ 9.230000000e-08 V_hig
+ 9.230100000e-08 V_hig
+ 9.240000000e-08 V_hig
+ 9.240100000e-08 V_hig
+ 9.250000000e-08 V_hig
+ 9.250100000e-08 V_hig
+ 9.260000000e-08 V_hig
+ 9.260100000e-08 V_hig
+ 9.270000000e-08 V_hig
+ 9.270100000e-08 V_hig
+ 9.280000000e-08 V_hig
+ 9.280100000e-08 V_hig
+ 9.290000000e-08 V_hig
+ 9.290100000e-08 V_low
+ 9.300000000e-08 V_low
+ 9.300100000e-08 V_low
+ 9.310000000e-08 V_low
+ 9.310100000e-08 V_low
+ 9.320000000e-08 V_low
+ 9.320100000e-08 V_low
+ 9.330000000e-08 V_low
+ 9.330100000e-08 V_low
+ 9.340000000e-08 V_low
+ 9.340100000e-08 V_low
+ 9.350000000e-08 V_low
+ 9.350100000e-08 V_low
+ 9.360000000e-08 V_low
+ 9.360100000e-08 V_low
+ 9.370000000e-08 V_low
+ 9.370100000e-08 V_low
+ 9.380000000e-08 V_low
+ 9.380100000e-08 V_low
+ 9.390000000e-08 V_low
+ 9.390100000e-08 V_hig
+ 9.400000000e-08 V_hig
+ 9.400100000e-08 V_hig
+ 9.410000000e-08 V_hig
+ 9.410100000e-08 V_hig
+ 9.420000000e-08 V_hig
+ 9.420100000e-08 V_hig
+ 9.430000000e-08 V_hig
+ 9.430100000e-08 V_hig
+ 9.440000000e-08 V_hig
+ 9.440100000e-08 V_hig
+ 9.450000000e-08 V_hig
+ 9.450100000e-08 V_hig
+ 9.460000000e-08 V_hig
+ 9.460100000e-08 V_hig
+ 9.470000000e-08 V_hig
+ 9.470100000e-08 V_hig
+ 9.480000000e-08 V_hig
+ 9.480100000e-08 V_hig
+ 9.490000000e-08 V_hig
+ 9.490100000e-08 V_hig
+ 9.500000000e-08 V_hig
+ 9.500100000e-08 V_hig
+ 9.510000000e-08 V_hig
+ 9.510100000e-08 V_hig
+ 9.520000000e-08 V_hig
+ 9.520100000e-08 V_hig
+ 9.530000000e-08 V_hig
+ 9.530100000e-08 V_hig
+ 9.540000000e-08 V_hig
+ 9.540100000e-08 V_hig
+ 9.550000000e-08 V_hig
+ 9.550100000e-08 V_hig
+ 9.560000000e-08 V_hig
+ 9.560100000e-08 V_hig
+ 9.570000000e-08 V_hig
+ 9.570100000e-08 V_hig
+ 9.580000000e-08 V_hig
+ 9.580100000e-08 V_hig
+ 9.590000000e-08 V_hig
+ 9.590100000e-08 V_low
+ 9.600000000e-08 V_low
+ 9.600100000e-08 V_low
+ 9.610000000e-08 V_low
+ 9.610100000e-08 V_low
+ 9.620000000e-08 V_low
+ 9.620100000e-08 V_low
+ 9.630000000e-08 V_low
+ 9.630100000e-08 V_low
+ 9.640000000e-08 V_low
+ 9.640100000e-08 V_low
+ 9.650000000e-08 V_low
+ 9.650100000e-08 V_low
+ 9.660000000e-08 V_low
+ 9.660100000e-08 V_low
+ 9.670000000e-08 V_low
+ 9.670100000e-08 V_low
+ 9.680000000e-08 V_low
+ 9.680100000e-08 V_low
+ 9.690000000e-08 V_low
+ 9.690100000e-08 V_low
+ 9.700000000e-08 V_low
+ 9.700100000e-08 V_low
+ 9.710000000e-08 V_low
+ 9.710100000e-08 V_low
+ 9.720000000e-08 V_low
+ 9.720100000e-08 V_low
+ 9.730000000e-08 V_low
+ 9.730100000e-08 V_low
+ 9.740000000e-08 V_low
+ 9.740100000e-08 V_low
+ 9.750000000e-08 V_low
+ 9.750100000e-08 V_low
+ 9.760000000e-08 V_low
+ 9.760100000e-08 V_low
+ 9.770000000e-08 V_low
+ 9.770100000e-08 V_low
+ 9.780000000e-08 V_low
+ 9.780100000e-08 V_low
+ 9.790000000e-08 V_low
+ 9.790100000e-08 V_hig
+ 9.800000000e-08 V_hig
+ 9.800100000e-08 V_hig
+ 9.810000000e-08 V_hig
+ 9.810100000e-08 V_hig
+ 9.820000000e-08 V_hig
+ 9.820100000e-08 V_hig
+ 9.830000000e-08 V_hig
+ 9.830100000e-08 V_hig
+ 9.840000000e-08 V_hig
+ 9.840100000e-08 V_hig
+ 9.850000000e-08 V_hig
+ 9.850100000e-08 V_hig
+ 9.860000000e-08 V_hig
+ 9.860100000e-08 V_hig
+ 9.870000000e-08 V_hig
+ 9.870100000e-08 V_hig
+ 9.880000000e-08 V_hig
+ 9.880100000e-08 V_hig
+ 9.890000000e-08 V_hig
+ 9.890100000e-08 V_hig
+ 9.900000000e-08 V_hig
+ 9.900100000e-08 V_hig
+ 9.910000000e-08 V_hig
+ 9.910100000e-08 V_hig
+ 9.920000000e-08 V_hig
+ 9.920100000e-08 V_hig
+ 9.930000000e-08 V_hig
+ 9.930100000e-08 V_hig
+ 9.940000000e-08 V_hig
+ 9.940100000e-08 V_hig
+ 9.950000000e-08 V_hig
+ 9.950100000e-08 V_hig
+ 9.960000000e-08 V_hig
+ 9.960100000e-08 V_hig
+ 9.970000000e-08 V_hig
+ 9.970100000e-08 V_hig
+ 9.980000000e-08 V_hig
+ 9.980100000e-08 V_hig
+ 9.990000000e-08 V_hig
+ 9.990100000e-08 V_hig
+ 1.000000000e-07 V_hig
+ 1.000010000e-07 V_hig
+ 1.001000000e-07 V_hig
+ 1.001010000e-07 V_hig
+ 1.002000000e-07 V_hig
+ 1.002010000e-07 V_hig
+ 1.003000000e-07 V_hig
+ 1.003010000e-07 V_hig
+ 1.004000000e-07 V_hig
+ 1.004010000e-07 V_hig
+ 1.005000000e-07 V_hig
+ 1.005010000e-07 V_hig
+ 1.006000000e-07 V_hig
+ 1.006010000e-07 V_hig
+ 1.007000000e-07 V_hig
+ 1.007010000e-07 V_hig
+ 1.008000000e-07 V_hig
+ 1.008010000e-07 V_hig
+ 1.009000000e-07 V_hig
+ 1.009010000e-07 V_hig
+ 1.010000000e-07 V_hig
+ 1.010010000e-07 V_hig
+ 1.011000000e-07 V_hig
+ 1.011010000e-07 V_hig
+ 1.012000000e-07 V_hig
+ 1.012010000e-07 V_hig
+ 1.013000000e-07 V_hig
+ 1.013010000e-07 V_hig
+ 1.014000000e-07 V_hig
+ 1.014010000e-07 V_hig
+ 1.015000000e-07 V_hig
+ 1.015010000e-07 V_hig
+ 1.016000000e-07 V_hig
+ 1.016010000e-07 V_hig
+ 1.017000000e-07 V_hig
+ 1.017010000e-07 V_hig
+ 1.018000000e-07 V_hig
+ 1.018010000e-07 V_hig
+ 1.019000000e-07 V_hig
+ 1.019010000e-07 V_hig
+ 1.020000000e-07 V_hig
+ 1.020010000e-07 V_hig
+ 1.021000000e-07 V_hig
+ 1.021010000e-07 V_hig
+ 1.022000000e-07 V_hig
+ 1.022010000e-07 V_hig
+ 1.023000000e-07 V_hig
+ 1.023010000e-07 V_hig
+ 1.024000000e-07 V_hig
+ 1.024010000e-07 V_hig
+ 1.025000000e-07 V_hig
+ 1.025010000e-07 V_hig
+ 1.026000000e-07 V_hig
+ 1.026010000e-07 V_hig
+ 1.027000000e-07 V_hig
+ 1.027010000e-07 V_hig
+ 1.028000000e-07 V_hig
+ 1.028010000e-07 V_hig
+ 1.029000000e-07 V_hig
+ 1.029010000e-07 V_low
+ 1.030000000e-07 V_low
+ 1.030010000e-07 V_low
+ 1.031000000e-07 V_low
+ 1.031010000e-07 V_low
+ 1.032000000e-07 V_low
+ 1.032010000e-07 V_low
+ 1.033000000e-07 V_low
+ 1.033010000e-07 V_low
+ 1.034000000e-07 V_low
+ 1.034010000e-07 V_low
+ 1.035000000e-07 V_low
+ 1.035010000e-07 V_low
+ 1.036000000e-07 V_low
+ 1.036010000e-07 V_low
+ 1.037000000e-07 V_low
+ 1.037010000e-07 V_low
+ 1.038000000e-07 V_low
+ 1.038010000e-07 V_low
+ 1.039000000e-07 V_low
+ 1.039010000e-07 V_hig
+ 1.040000000e-07 V_hig
+ 1.040010000e-07 V_hig
+ 1.041000000e-07 V_hig
+ 1.041010000e-07 V_hig
+ 1.042000000e-07 V_hig
+ 1.042010000e-07 V_hig
+ 1.043000000e-07 V_hig
+ 1.043010000e-07 V_hig
+ 1.044000000e-07 V_hig
+ 1.044010000e-07 V_hig
+ 1.045000000e-07 V_hig
+ 1.045010000e-07 V_hig
+ 1.046000000e-07 V_hig
+ 1.046010000e-07 V_hig
+ 1.047000000e-07 V_hig
+ 1.047010000e-07 V_hig
+ 1.048000000e-07 V_hig
+ 1.048010000e-07 V_hig
+ 1.049000000e-07 V_hig
+ 1.049010000e-07 V_hig
+ 1.050000000e-07 V_hig
+ 1.050010000e-07 V_hig
+ 1.051000000e-07 V_hig
+ 1.051010000e-07 V_hig
+ 1.052000000e-07 V_hig
+ 1.052010000e-07 V_hig
+ 1.053000000e-07 V_hig
+ 1.053010000e-07 V_hig
+ 1.054000000e-07 V_hig
+ 1.054010000e-07 V_hig
+ 1.055000000e-07 V_hig
+ 1.055010000e-07 V_hig
+ 1.056000000e-07 V_hig
+ 1.056010000e-07 V_hig
+ 1.057000000e-07 V_hig
+ 1.057010000e-07 V_hig
+ 1.058000000e-07 V_hig
+ 1.058010000e-07 V_hig
+ 1.059000000e-07 V_hig
+ 1.059010000e-07 V_hig
+ 1.060000000e-07 V_hig
+ 1.060010000e-07 V_hig
+ 1.061000000e-07 V_hig
+ 1.061010000e-07 V_hig
+ 1.062000000e-07 V_hig
+ 1.062010000e-07 V_hig
+ 1.063000000e-07 V_hig
+ 1.063010000e-07 V_hig
+ 1.064000000e-07 V_hig
+ 1.064010000e-07 V_hig
+ 1.065000000e-07 V_hig
+ 1.065010000e-07 V_hig
+ 1.066000000e-07 V_hig
+ 1.066010000e-07 V_hig
+ 1.067000000e-07 V_hig
+ 1.067010000e-07 V_hig
+ 1.068000000e-07 V_hig
+ 1.068010000e-07 V_hig
+ 1.069000000e-07 V_hig
+ 1.069010000e-07 V_hig
+ 1.070000000e-07 V_hig
+ 1.070010000e-07 V_hig
+ 1.071000000e-07 V_hig
+ 1.071010000e-07 V_hig
+ 1.072000000e-07 V_hig
+ 1.072010000e-07 V_hig
+ 1.073000000e-07 V_hig
+ 1.073010000e-07 V_hig
+ 1.074000000e-07 V_hig
+ 1.074010000e-07 V_hig
+ 1.075000000e-07 V_hig
+ 1.075010000e-07 V_hig
+ 1.076000000e-07 V_hig
+ 1.076010000e-07 V_hig
+ 1.077000000e-07 V_hig
+ 1.077010000e-07 V_hig
+ 1.078000000e-07 V_hig
+ 1.078010000e-07 V_hig
+ 1.079000000e-07 V_hig
+ 1.079010000e-07 V_low
+ 1.080000000e-07 V_low
+ 1.080010000e-07 V_low
+ 1.081000000e-07 V_low
+ 1.081010000e-07 V_low
+ 1.082000000e-07 V_low
+ 1.082010000e-07 V_low
+ 1.083000000e-07 V_low
+ 1.083010000e-07 V_low
+ 1.084000000e-07 V_low
+ 1.084010000e-07 V_low
+ 1.085000000e-07 V_low
+ 1.085010000e-07 V_low
+ 1.086000000e-07 V_low
+ 1.086010000e-07 V_low
+ 1.087000000e-07 V_low
+ 1.087010000e-07 V_low
+ 1.088000000e-07 V_low
+ 1.088010000e-07 V_low
+ 1.089000000e-07 V_low
+ 1.089010000e-07 V_low
+ 1.090000000e-07 V_low
+ 1.090010000e-07 V_low
+ 1.091000000e-07 V_low
+ 1.091010000e-07 V_low
+ 1.092000000e-07 V_low
+ 1.092010000e-07 V_low
+ 1.093000000e-07 V_low
+ 1.093010000e-07 V_low
+ 1.094000000e-07 V_low
+ 1.094010000e-07 V_low
+ 1.095000000e-07 V_low
+ 1.095010000e-07 V_low
+ 1.096000000e-07 V_low
+ 1.096010000e-07 V_low
+ 1.097000000e-07 V_low
+ 1.097010000e-07 V_low
+ 1.098000000e-07 V_low
+ 1.098010000e-07 V_low
+ 1.099000000e-07 V_low
+ 1.099010000e-07 V_low
+ 1.100000000e-07 V_low
+ 1.100010000e-07 V_low
+ 1.101000000e-07 V_low
+ 1.101010000e-07 V_low
+ 1.102000000e-07 V_low
+ 1.102010000e-07 V_low
+ 1.103000000e-07 V_low
+ 1.103010000e-07 V_low
+ 1.104000000e-07 V_low
+ 1.104010000e-07 V_low
+ 1.105000000e-07 V_low
+ 1.105010000e-07 V_low
+ 1.106000000e-07 V_low
+ 1.106010000e-07 V_low
+ 1.107000000e-07 V_low
+ 1.107010000e-07 V_low
+ 1.108000000e-07 V_low
+ 1.108010000e-07 V_low
+ 1.109000000e-07 V_low
+ 1.109010000e-07 V_low
+ 1.110000000e-07 V_low
+ 1.110010000e-07 V_low
+ 1.111000000e-07 V_low
+ 1.111010000e-07 V_low
+ 1.112000000e-07 V_low
+ 1.112010000e-07 V_low
+ 1.113000000e-07 V_low
+ 1.113010000e-07 V_low
+ 1.114000000e-07 V_low
+ 1.114010000e-07 V_low
+ 1.115000000e-07 V_low
+ 1.115010000e-07 V_low
+ 1.116000000e-07 V_low
+ 1.116010000e-07 V_low
+ 1.117000000e-07 V_low
+ 1.117010000e-07 V_low
+ 1.118000000e-07 V_low
+ 1.118010000e-07 V_low
+ 1.119000000e-07 V_low
+ 1.119010000e-07 V_hig
+ 1.120000000e-07 V_hig
+ 1.120010000e-07 V_hig
+ 1.121000000e-07 V_hig
+ 1.121010000e-07 V_hig
+ 1.122000000e-07 V_hig
+ 1.122010000e-07 V_hig
+ 1.123000000e-07 V_hig
+ 1.123010000e-07 V_hig
+ 1.124000000e-07 V_hig
+ 1.124010000e-07 V_hig
+ 1.125000000e-07 V_hig
+ 1.125010000e-07 V_hig
+ 1.126000000e-07 V_hig
+ 1.126010000e-07 V_hig
+ 1.127000000e-07 V_hig
+ 1.127010000e-07 V_hig
+ 1.128000000e-07 V_hig
+ 1.128010000e-07 V_hig
+ 1.129000000e-07 V_hig
+ 1.129010000e-07 V_low
+ 1.130000000e-07 V_low
+ 1.130010000e-07 V_low
+ 1.131000000e-07 V_low
+ 1.131010000e-07 V_low
+ 1.132000000e-07 V_low
+ 1.132010000e-07 V_low
+ 1.133000000e-07 V_low
+ 1.133010000e-07 V_low
+ 1.134000000e-07 V_low
+ 1.134010000e-07 V_low
+ 1.135000000e-07 V_low
+ 1.135010000e-07 V_low
+ 1.136000000e-07 V_low
+ 1.136010000e-07 V_low
+ 1.137000000e-07 V_low
+ 1.137010000e-07 V_low
+ 1.138000000e-07 V_low
+ 1.138010000e-07 V_low
+ 1.139000000e-07 V_low
+ 1.139010000e-07 V_low
+ 1.140000000e-07 V_low
+ 1.140010000e-07 V_low
+ 1.141000000e-07 V_low
+ 1.141010000e-07 V_low
+ 1.142000000e-07 V_low
+ 1.142010000e-07 V_low
+ 1.143000000e-07 V_low
+ 1.143010000e-07 V_low
+ 1.144000000e-07 V_low
+ 1.144010000e-07 V_low
+ 1.145000000e-07 V_low
+ 1.145010000e-07 V_low
+ 1.146000000e-07 V_low
+ 1.146010000e-07 V_low
+ 1.147000000e-07 V_low
+ 1.147010000e-07 V_low
+ 1.148000000e-07 V_low
+ 1.148010000e-07 V_low
+ 1.149000000e-07 V_low
+ 1.149010000e-07 V_hig
+ 1.150000000e-07 V_hig
+ 1.150010000e-07 V_hig
+ 1.151000000e-07 V_hig
+ 1.151010000e-07 V_hig
+ 1.152000000e-07 V_hig
+ 1.152010000e-07 V_hig
+ 1.153000000e-07 V_hig
+ 1.153010000e-07 V_hig
+ 1.154000000e-07 V_hig
+ 1.154010000e-07 V_hig
+ 1.155000000e-07 V_hig
+ 1.155010000e-07 V_hig
+ 1.156000000e-07 V_hig
+ 1.156010000e-07 V_hig
+ 1.157000000e-07 V_hig
+ 1.157010000e-07 V_hig
+ 1.158000000e-07 V_hig
+ 1.158010000e-07 V_hig
+ 1.159000000e-07 V_hig
+ 1.159010000e-07 V_hig
+ 1.160000000e-07 V_hig
+ 1.160010000e-07 V_hig
+ 1.161000000e-07 V_hig
+ 1.161010000e-07 V_hig
+ 1.162000000e-07 V_hig
+ 1.162010000e-07 V_hig
+ 1.163000000e-07 V_hig
+ 1.163010000e-07 V_hig
+ 1.164000000e-07 V_hig
+ 1.164010000e-07 V_hig
+ 1.165000000e-07 V_hig
+ 1.165010000e-07 V_hig
+ 1.166000000e-07 V_hig
+ 1.166010000e-07 V_hig
+ 1.167000000e-07 V_hig
+ 1.167010000e-07 V_hig
+ 1.168000000e-07 V_hig
+ 1.168010000e-07 V_hig
+ 1.169000000e-07 V_hig
+ 1.169010000e-07 V_hig
+ 1.170000000e-07 V_hig
+ 1.170010000e-07 V_hig
+ 1.171000000e-07 V_hig
+ 1.171010000e-07 V_hig
+ 1.172000000e-07 V_hig
+ 1.172010000e-07 V_hig
+ 1.173000000e-07 V_hig
+ 1.173010000e-07 V_hig
+ 1.174000000e-07 V_hig
+ 1.174010000e-07 V_hig
+ 1.175000000e-07 V_hig
+ 1.175010000e-07 V_hig
+ 1.176000000e-07 V_hig
+ 1.176010000e-07 V_hig
+ 1.177000000e-07 V_hig
+ 1.177010000e-07 V_hig
+ 1.178000000e-07 V_hig
+ 1.178010000e-07 V_hig
+ 1.179000000e-07 V_hig
+ 1.179010000e-07 V_low
+ 1.180000000e-07 V_low
+ 1.180010000e-07 V_low
+ 1.181000000e-07 V_low
+ 1.181010000e-07 V_low
+ 1.182000000e-07 V_low
+ 1.182010000e-07 V_low
+ 1.183000000e-07 V_low
+ 1.183010000e-07 V_low
+ 1.184000000e-07 V_low
+ 1.184010000e-07 V_low
+ 1.185000000e-07 V_low
+ 1.185010000e-07 V_low
+ 1.186000000e-07 V_low
+ 1.186010000e-07 V_low
+ 1.187000000e-07 V_low
+ 1.187010000e-07 V_low
+ 1.188000000e-07 V_low
+ 1.188010000e-07 V_low
+ 1.189000000e-07 V_low
+ 1.189010000e-07 V_low
+ 1.190000000e-07 V_low
+ 1.190010000e-07 V_low
+ 1.191000000e-07 V_low
+ 1.191010000e-07 V_low
+ 1.192000000e-07 V_low
+ 1.192010000e-07 V_low
+ 1.193000000e-07 V_low
+ 1.193010000e-07 V_low
+ 1.194000000e-07 V_low
+ 1.194010000e-07 V_low
+ 1.195000000e-07 V_low
+ 1.195010000e-07 V_low
+ 1.196000000e-07 V_low
+ 1.196010000e-07 V_low
+ 1.197000000e-07 V_low
+ 1.197010000e-07 V_low
+ 1.198000000e-07 V_low
+ 1.198010000e-07 V_low
+ 1.199000000e-07 V_low
+ 1.199010000e-07 V_low
+ 1.200000000e-07 V_low
+ 1.200010000e-07 V_low
+ 1.201000000e-07 V_low
+ 1.201010000e-07 V_low
+ 1.202000000e-07 V_low
+ 1.202010000e-07 V_low
+ 1.203000000e-07 V_low
+ 1.203010000e-07 V_low
+ 1.204000000e-07 V_low
+ 1.204010000e-07 V_low
+ 1.205000000e-07 V_low
+ 1.205010000e-07 V_low
+ 1.206000000e-07 V_low
+ 1.206010000e-07 V_low
+ 1.207000000e-07 V_low
+ 1.207010000e-07 V_low
+ 1.208000000e-07 V_low
+ 1.208010000e-07 V_low
+ 1.209000000e-07 V_low
+ 1.209010000e-07 V_hig
+ 1.210000000e-07 V_hig
+ 1.210010000e-07 V_hig
+ 1.211000000e-07 V_hig
+ 1.211010000e-07 V_hig
+ 1.212000000e-07 V_hig
+ 1.212010000e-07 V_hig
+ 1.213000000e-07 V_hig
+ 1.213010000e-07 V_hig
+ 1.214000000e-07 V_hig
+ 1.214010000e-07 V_hig
+ 1.215000000e-07 V_hig
+ 1.215010000e-07 V_hig
+ 1.216000000e-07 V_hig
+ 1.216010000e-07 V_hig
+ 1.217000000e-07 V_hig
+ 1.217010000e-07 V_hig
+ 1.218000000e-07 V_hig
+ 1.218010000e-07 V_hig
+ 1.219000000e-07 V_hig
+ 1.219010000e-07 V_hig
+ 1.220000000e-07 V_hig
+ 1.220010000e-07 V_hig
+ 1.221000000e-07 V_hig
+ 1.221010000e-07 V_hig
+ 1.222000000e-07 V_hig
+ 1.222010000e-07 V_hig
+ 1.223000000e-07 V_hig
+ 1.223010000e-07 V_hig
+ 1.224000000e-07 V_hig
+ 1.224010000e-07 V_hig
+ 1.225000000e-07 V_hig
+ 1.225010000e-07 V_hig
+ 1.226000000e-07 V_hig
+ 1.226010000e-07 V_hig
+ 1.227000000e-07 V_hig
+ 1.227010000e-07 V_hig
+ 1.228000000e-07 V_hig
+ 1.228010000e-07 V_hig
+ 1.229000000e-07 V_hig
+ 1.229010000e-07 V_hig
+ 1.230000000e-07 V_hig
+ 1.230010000e-07 V_hig
+ 1.231000000e-07 V_hig
+ 1.231010000e-07 V_hig
+ 1.232000000e-07 V_hig
+ 1.232010000e-07 V_hig
+ 1.233000000e-07 V_hig
+ 1.233010000e-07 V_hig
+ 1.234000000e-07 V_hig
+ 1.234010000e-07 V_hig
+ 1.235000000e-07 V_hig
+ 1.235010000e-07 V_hig
+ 1.236000000e-07 V_hig
+ 1.236010000e-07 V_hig
+ 1.237000000e-07 V_hig
+ 1.237010000e-07 V_hig
+ 1.238000000e-07 V_hig
+ 1.238010000e-07 V_hig
+ 1.239000000e-07 V_hig
+ 1.239010000e-07 V_low
+ 1.240000000e-07 V_low
+ 1.240010000e-07 V_low
+ 1.241000000e-07 V_low
+ 1.241010000e-07 V_low
+ 1.242000000e-07 V_low
+ 1.242010000e-07 V_low
+ 1.243000000e-07 V_low
+ 1.243010000e-07 V_low
+ 1.244000000e-07 V_low
+ 1.244010000e-07 V_low
+ 1.245000000e-07 V_low
+ 1.245010000e-07 V_low
+ 1.246000000e-07 V_low
+ 1.246010000e-07 V_low
+ 1.247000000e-07 V_low
+ 1.247010000e-07 V_low
+ 1.248000000e-07 V_low
+ 1.248010000e-07 V_low
+ 1.249000000e-07 V_low
+ 1.249010000e-07 V_hig
+ 1.250000000e-07 V_hig
+ 1.250010000e-07 V_hig
+ 1.251000000e-07 V_hig
+ 1.251010000e-07 V_hig
+ 1.252000000e-07 V_hig
+ 1.252010000e-07 V_hig
+ 1.253000000e-07 V_hig
+ 1.253010000e-07 V_hig
+ 1.254000000e-07 V_hig
+ 1.254010000e-07 V_hig
+ 1.255000000e-07 V_hig
+ 1.255010000e-07 V_hig
+ 1.256000000e-07 V_hig
+ 1.256010000e-07 V_hig
+ 1.257000000e-07 V_hig
+ 1.257010000e-07 V_hig
+ 1.258000000e-07 V_hig
+ 1.258010000e-07 V_hig
+ 1.259000000e-07 V_hig
+ 1.259010000e-07 V_low
+ 1.260000000e-07 V_low
+ 1.260010000e-07 V_low
+ 1.261000000e-07 V_low
+ 1.261010000e-07 V_low
+ 1.262000000e-07 V_low
+ 1.262010000e-07 V_low
+ 1.263000000e-07 V_low
+ 1.263010000e-07 V_low
+ 1.264000000e-07 V_low
+ 1.264010000e-07 V_low
+ 1.265000000e-07 V_low
+ 1.265010000e-07 V_low
+ 1.266000000e-07 V_low
+ 1.266010000e-07 V_low
+ 1.267000000e-07 V_low
+ 1.267010000e-07 V_low
+ 1.268000000e-07 V_low
+ 1.268010000e-07 V_low
+ 1.269000000e-07 V_low
+ 1.269010000e-07 V_low
+ 1.270000000e-07 V_low
+ 1.270010000e-07 V_low
+ 1.271000000e-07 V_low
+ 1.271010000e-07 V_low
+ 1.272000000e-07 V_low
+ 1.272010000e-07 V_low
+ 1.273000000e-07 V_low
+ 1.273010000e-07 V_low
+ 1.274000000e-07 V_low
+ 1.274010000e-07 V_low
+ 1.275000000e-07 V_low
+ 1.275010000e-07 V_low
+ 1.276000000e-07 V_low
+ 1.276010000e-07 V_low
+ 1.277000000e-07 V_low
+ 1.277010000e-07 V_low
+ 1.278000000e-07 V_low
+ 1.278010000e-07 V_low
+ 1.279000000e-07 V_low
+ 1.279010000e-07 V_low
+ 1.280000000e-07 V_low
+ 1.280010000e-07 V_low
+ 1.281000000e-07 V_low
+ 1.281010000e-07 V_low
+ 1.282000000e-07 V_low
+ 1.282010000e-07 V_low
+ 1.283000000e-07 V_low
+ 1.283010000e-07 V_low
+ 1.284000000e-07 V_low
+ 1.284010000e-07 V_low
+ 1.285000000e-07 V_low
+ 1.285010000e-07 V_low
+ 1.286000000e-07 V_low
+ 1.286010000e-07 V_low
+ 1.287000000e-07 V_low
+ 1.287010000e-07 V_low
+ 1.288000000e-07 V_low
+ 1.288010000e-07 V_low
+ 1.289000000e-07 V_low
+ 1.289010000e-07 V_low
+ 1.290000000e-07 V_low
+ 1.290010000e-07 V_low
+ 1.291000000e-07 V_low
+ 1.291010000e-07 V_low
+ 1.292000000e-07 V_low
+ 1.292010000e-07 V_low
+ 1.293000000e-07 V_low
+ 1.293010000e-07 V_low
+ 1.294000000e-07 V_low
+ 1.294010000e-07 V_low
+ 1.295000000e-07 V_low
+ 1.295010000e-07 V_low
+ 1.296000000e-07 V_low
+ 1.296010000e-07 V_low
+ 1.297000000e-07 V_low
+ 1.297010000e-07 V_low
+ 1.298000000e-07 V_low
+ 1.298010000e-07 V_low
+ 1.299000000e-07 V_low
+ 1.299010000e-07 V_hig
+ 1.300000000e-07 V_hig
+ 1.300010000e-07 V_hig
+ 1.301000000e-07 V_hig
+ 1.301010000e-07 V_hig
+ 1.302000000e-07 V_hig
+ 1.302010000e-07 V_hig
+ 1.303000000e-07 V_hig
+ 1.303010000e-07 V_hig
+ 1.304000000e-07 V_hig
+ 1.304010000e-07 V_hig
+ 1.305000000e-07 V_hig
+ 1.305010000e-07 V_hig
+ 1.306000000e-07 V_hig
+ 1.306010000e-07 V_hig
+ 1.307000000e-07 V_hig
+ 1.307010000e-07 V_hig
+ 1.308000000e-07 V_hig
+ 1.308010000e-07 V_hig
+ 1.309000000e-07 V_hig
+ 1.309010000e-07 V_hig
+ 1.310000000e-07 V_hig
+ 1.310010000e-07 V_hig
+ 1.311000000e-07 V_hig
+ 1.311010000e-07 V_hig
+ 1.312000000e-07 V_hig
+ 1.312010000e-07 V_hig
+ 1.313000000e-07 V_hig
+ 1.313010000e-07 V_hig
+ 1.314000000e-07 V_hig
+ 1.314010000e-07 V_hig
+ 1.315000000e-07 V_hig
+ 1.315010000e-07 V_hig
+ 1.316000000e-07 V_hig
+ 1.316010000e-07 V_hig
+ 1.317000000e-07 V_hig
+ 1.317010000e-07 V_hig
+ 1.318000000e-07 V_hig
+ 1.318010000e-07 V_hig
+ 1.319000000e-07 V_hig
+ 1.319010000e-07 V_hig
+ 1.320000000e-07 V_hig
+ 1.320010000e-07 V_hig
+ 1.321000000e-07 V_hig
+ 1.321010000e-07 V_hig
+ 1.322000000e-07 V_hig
+ 1.322010000e-07 V_hig
+ 1.323000000e-07 V_hig
+ 1.323010000e-07 V_hig
+ 1.324000000e-07 V_hig
+ 1.324010000e-07 V_hig
+ 1.325000000e-07 V_hig
+ 1.325010000e-07 V_hig
+ 1.326000000e-07 V_hig
+ 1.326010000e-07 V_hig
+ 1.327000000e-07 V_hig
+ 1.327010000e-07 V_hig
+ 1.328000000e-07 V_hig
+ 1.328010000e-07 V_hig
+ 1.329000000e-07 V_hig
+ 1.329010000e-07 V_low
+ 1.330000000e-07 V_low
+ 1.330010000e-07 V_low
+ 1.331000000e-07 V_low
+ 1.331010000e-07 V_low
+ 1.332000000e-07 V_low
+ 1.332010000e-07 V_low
+ 1.333000000e-07 V_low
+ 1.333010000e-07 V_low
+ 1.334000000e-07 V_low
+ 1.334010000e-07 V_low
+ 1.335000000e-07 V_low
+ 1.335010000e-07 V_low
+ 1.336000000e-07 V_low
+ 1.336010000e-07 V_low
+ 1.337000000e-07 V_low
+ 1.337010000e-07 V_low
+ 1.338000000e-07 V_low
+ 1.338010000e-07 V_low
+ 1.339000000e-07 V_low
+ 1.339010000e-07 V_hig
+ 1.340000000e-07 V_hig
+ 1.340010000e-07 V_hig
+ 1.341000000e-07 V_hig
+ 1.341010000e-07 V_hig
+ 1.342000000e-07 V_hig
+ 1.342010000e-07 V_hig
+ 1.343000000e-07 V_hig
+ 1.343010000e-07 V_hig
+ 1.344000000e-07 V_hig
+ 1.344010000e-07 V_hig
+ 1.345000000e-07 V_hig
+ 1.345010000e-07 V_hig
+ 1.346000000e-07 V_hig
+ 1.346010000e-07 V_hig
+ 1.347000000e-07 V_hig
+ 1.347010000e-07 V_hig
+ 1.348000000e-07 V_hig
+ 1.348010000e-07 V_hig
+ 1.349000000e-07 V_hig
+ 1.349010000e-07 V_low
+ 1.350000000e-07 V_low
+ 1.350010000e-07 V_low
+ 1.351000000e-07 V_low
+ 1.351010000e-07 V_low
+ 1.352000000e-07 V_low
+ 1.352010000e-07 V_low
+ 1.353000000e-07 V_low
+ 1.353010000e-07 V_low
+ 1.354000000e-07 V_low
+ 1.354010000e-07 V_low
+ 1.355000000e-07 V_low
+ 1.355010000e-07 V_low
+ 1.356000000e-07 V_low
+ 1.356010000e-07 V_low
+ 1.357000000e-07 V_low
+ 1.357010000e-07 V_low
+ 1.358000000e-07 V_low
+ 1.358010000e-07 V_low
+ 1.359000000e-07 V_low
+ 1.359010000e-07 V_hig
+ 1.360000000e-07 V_hig
+ 1.360010000e-07 V_hig
+ 1.361000000e-07 V_hig
+ 1.361010000e-07 V_hig
+ 1.362000000e-07 V_hig
+ 1.362010000e-07 V_hig
+ 1.363000000e-07 V_hig
+ 1.363010000e-07 V_hig
+ 1.364000000e-07 V_hig
+ 1.364010000e-07 V_hig
+ 1.365000000e-07 V_hig
+ 1.365010000e-07 V_hig
+ 1.366000000e-07 V_hig
+ 1.366010000e-07 V_hig
+ 1.367000000e-07 V_hig
+ 1.367010000e-07 V_hig
+ 1.368000000e-07 V_hig
+ 1.368010000e-07 V_hig
+ 1.369000000e-07 V_hig
+ 1.369010000e-07 V_low
+ 1.370000000e-07 V_low
+ 1.370010000e-07 V_low
+ 1.371000000e-07 V_low
+ 1.371010000e-07 V_low
+ 1.372000000e-07 V_low
+ 1.372010000e-07 V_low
+ 1.373000000e-07 V_low
+ 1.373010000e-07 V_low
+ 1.374000000e-07 V_low
+ 1.374010000e-07 V_low
+ 1.375000000e-07 V_low
+ 1.375010000e-07 V_low
+ 1.376000000e-07 V_low
+ 1.376010000e-07 V_low
+ 1.377000000e-07 V_low
+ 1.377010000e-07 V_low
+ 1.378000000e-07 V_low
+ 1.378010000e-07 V_low
+ 1.379000000e-07 V_low
+ 1.379010000e-07 V_hig
+ 1.380000000e-07 V_hig
+ 1.380010000e-07 V_hig
+ 1.381000000e-07 V_hig
+ 1.381010000e-07 V_hig
+ 1.382000000e-07 V_hig
+ 1.382010000e-07 V_hig
+ 1.383000000e-07 V_hig
+ 1.383010000e-07 V_hig
+ 1.384000000e-07 V_hig
+ 1.384010000e-07 V_hig
+ 1.385000000e-07 V_hig
+ 1.385010000e-07 V_hig
+ 1.386000000e-07 V_hig
+ 1.386010000e-07 V_hig
+ 1.387000000e-07 V_hig
+ 1.387010000e-07 V_hig
+ 1.388000000e-07 V_hig
+ 1.388010000e-07 V_hig
+ 1.389000000e-07 V_hig
+ 1.389010000e-07 V_hig
+ 1.390000000e-07 V_hig
+ 1.390010000e-07 V_hig
+ 1.391000000e-07 V_hig
+ 1.391010000e-07 V_hig
+ 1.392000000e-07 V_hig
+ 1.392010000e-07 V_hig
+ 1.393000000e-07 V_hig
+ 1.393010000e-07 V_hig
+ 1.394000000e-07 V_hig
+ 1.394010000e-07 V_hig
+ 1.395000000e-07 V_hig
+ 1.395010000e-07 V_hig
+ 1.396000000e-07 V_hig
+ 1.396010000e-07 V_hig
+ 1.397000000e-07 V_hig
+ 1.397010000e-07 V_hig
+ 1.398000000e-07 V_hig
+ 1.398010000e-07 V_hig
+ 1.399000000e-07 V_hig
+ 1.399010000e-07 V_hig
+ 1.400000000e-07 V_hig
+ 1.400010000e-07 V_hig
+ 1.401000000e-07 V_hig
+ 1.401010000e-07 V_hig
+ 1.402000000e-07 V_hig
+ 1.402010000e-07 V_hig
+ 1.403000000e-07 V_hig
+ 1.403010000e-07 V_hig
+ 1.404000000e-07 V_hig
+ 1.404010000e-07 V_hig
+ 1.405000000e-07 V_hig
+ 1.405010000e-07 V_hig
+ 1.406000000e-07 V_hig
+ 1.406010000e-07 V_hig
+ 1.407000000e-07 V_hig
+ 1.407010000e-07 V_hig
+ 1.408000000e-07 V_hig
+ 1.408010000e-07 V_hig
+ 1.409000000e-07 V_hig
+ 1.409010000e-07 V_low
+ 1.410000000e-07 V_low
+ 1.410010000e-07 V_low
+ 1.411000000e-07 V_low
+ 1.411010000e-07 V_low
+ 1.412000000e-07 V_low
+ 1.412010000e-07 V_low
+ 1.413000000e-07 V_low
+ 1.413010000e-07 V_low
+ 1.414000000e-07 V_low
+ 1.414010000e-07 V_low
+ 1.415000000e-07 V_low
+ 1.415010000e-07 V_low
+ 1.416000000e-07 V_low
+ 1.416010000e-07 V_low
+ 1.417000000e-07 V_low
+ 1.417010000e-07 V_low
+ 1.418000000e-07 V_low
+ 1.418010000e-07 V_low
+ 1.419000000e-07 V_low
+ 1.419010000e-07 V_low
+ 1.420000000e-07 V_low
+ 1.420010000e-07 V_low
+ 1.421000000e-07 V_low
+ 1.421010000e-07 V_low
+ 1.422000000e-07 V_low
+ 1.422010000e-07 V_low
+ 1.423000000e-07 V_low
+ 1.423010000e-07 V_low
+ 1.424000000e-07 V_low
+ 1.424010000e-07 V_low
+ 1.425000000e-07 V_low
+ 1.425010000e-07 V_low
+ 1.426000000e-07 V_low
+ 1.426010000e-07 V_low
+ 1.427000000e-07 V_low
+ 1.427010000e-07 V_low
+ 1.428000000e-07 V_low
+ 1.428010000e-07 V_low
+ 1.429000000e-07 V_low
+ 1.429010000e-07 V_hig
+ 1.430000000e-07 V_hig
+ 1.430010000e-07 V_hig
+ 1.431000000e-07 V_hig
+ 1.431010000e-07 V_hig
+ 1.432000000e-07 V_hig
+ 1.432010000e-07 V_hig
+ 1.433000000e-07 V_hig
+ 1.433010000e-07 V_hig
+ 1.434000000e-07 V_hig
+ 1.434010000e-07 V_hig
+ 1.435000000e-07 V_hig
+ 1.435010000e-07 V_hig
+ 1.436000000e-07 V_hig
+ 1.436010000e-07 V_hig
+ 1.437000000e-07 V_hig
+ 1.437010000e-07 V_hig
+ 1.438000000e-07 V_hig
+ 1.438010000e-07 V_hig
+ 1.439000000e-07 V_hig
+ 1.439010000e-07 V_low
+ 1.440000000e-07 V_low
+ 1.440010000e-07 V_low
+ 1.441000000e-07 V_low
+ 1.441010000e-07 V_low
+ 1.442000000e-07 V_low
+ 1.442010000e-07 V_low
+ 1.443000000e-07 V_low
+ 1.443010000e-07 V_low
+ 1.444000000e-07 V_low
+ 1.444010000e-07 V_low
+ 1.445000000e-07 V_low
+ 1.445010000e-07 V_low
+ 1.446000000e-07 V_low
+ 1.446010000e-07 V_low
+ 1.447000000e-07 V_low
+ 1.447010000e-07 V_low
+ 1.448000000e-07 V_low
+ 1.448010000e-07 V_low
+ 1.449000000e-07 V_low
+ 1.449010000e-07 V_hig
+ 1.450000000e-07 V_hig
+ 1.450010000e-07 V_hig
+ 1.451000000e-07 V_hig
+ 1.451010000e-07 V_hig
+ 1.452000000e-07 V_hig
+ 1.452010000e-07 V_hig
+ 1.453000000e-07 V_hig
+ 1.453010000e-07 V_hig
+ 1.454000000e-07 V_hig
+ 1.454010000e-07 V_hig
+ 1.455000000e-07 V_hig
+ 1.455010000e-07 V_hig
+ 1.456000000e-07 V_hig
+ 1.456010000e-07 V_hig
+ 1.457000000e-07 V_hig
+ 1.457010000e-07 V_hig
+ 1.458000000e-07 V_hig
+ 1.458010000e-07 V_hig
+ 1.459000000e-07 V_hig
+ 1.459010000e-07 V_hig
+ 1.460000000e-07 V_hig
+ 1.460010000e-07 V_hig
+ 1.461000000e-07 V_hig
+ 1.461010000e-07 V_hig
+ 1.462000000e-07 V_hig
+ 1.462010000e-07 V_hig
+ 1.463000000e-07 V_hig
+ 1.463010000e-07 V_hig
+ 1.464000000e-07 V_hig
+ 1.464010000e-07 V_hig
+ 1.465000000e-07 V_hig
+ 1.465010000e-07 V_hig
+ 1.466000000e-07 V_hig
+ 1.466010000e-07 V_hig
+ 1.467000000e-07 V_hig
+ 1.467010000e-07 V_hig
+ 1.468000000e-07 V_hig
+ 1.468010000e-07 V_hig
+ 1.469000000e-07 V_hig
+ 1.469010000e-07 V_low
+ 1.470000000e-07 V_low
+ 1.470010000e-07 V_low
+ 1.471000000e-07 V_low
+ 1.471010000e-07 V_low
+ 1.472000000e-07 V_low
+ 1.472010000e-07 V_low
+ 1.473000000e-07 V_low
+ 1.473010000e-07 V_low
+ 1.474000000e-07 V_low
+ 1.474010000e-07 V_low
+ 1.475000000e-07 V_low
+ 1.475010000e-07 V_low
+ 1.476000000e-07 V_low
+ 1.476010000e-07 V_low
+ 1.477000000e-07 V_low
+ 1.477010000e-07 V_low
+ 1.478000000e-07 V_low
+ 1.478010000e-07 V_low
+ 1.479000000e-07 V_low
+ 1.479010000e-07 V_low
+ 1.480000000e-07 V_low
+ 1.480010000e-07 V_low
+ 1.481000000e-07 V_low
+ 1.481010000e-07 V_low
+ 1.482000000e-07 V_low
+ 1.482010000e-07 V_low
+ 1.483000000e-07 V_low
+ 1.483010000e-07 V_low
+ 1.484000000e-07 V_low
+ 1.484010000e-07 V_low
+ 1.485000000e-07 V_low
+ 1.485010000e-07 V_low
+ 1.486000000e-07 V_low
+ 1.486010000e-07 V_low
+ 1.487000000e-07 V_low
+ 1.487010000e-07 V_low
+ 1.488000000e-07 V_low
+ 1.488010000e-07 V_low
+ 1.489000000e-07 V_low
+ 1.489010000e-07 V_low
+ 1.490000000e-07 V_low
+ 1.490010000e-07 V_low
+ 1.491000000e-07 V_low
+ 1.491010000e-07 V_low
+ 1.492000000e-07 V_low
+ 1.492010000e-07 V_low
+ 1.493000000e-07 V_low
+ 1.493010000e-07 V_low
+ 1.494000000e-07 V_low
+ 1.494010000e-07 V_low
+ 1.495000000e-07 V_low
+ 1.495010000e-07 V_low
+ 1.496000000e-07 V_low
+ 1.496010000e-07 V_low
+ 1.497000000e-07 V_low
+ 1.497010000e-07 V_low
+ 1.498000000e-07 V_low
+ 1.498010000e-07 V_low
+ 1.499000000e-07 V_low
+ 1.499010000e-07 V_low
+ 1.500000000e-07 V_low
+ 1.500010000e-07 V_low
+ 1.501000000e-07 V_low
+ 1.501010000e-07 V_low
+ 1.502000000e-07 V_low
+ 1.502010000e-07 V_low
+ 1.503000000e-07 V_low
+ 1.503010000e-07 V_low
+ 1.504000000e-07 V_low
+ 1.504010000e-07 V_low
+ 1.505000000e-07 V_low
+ 1.505010000e-07 V_low
+ 1.506000000e-07 V_low
+ 1.506010000e-07 V_low
+ 1.507000000e-07 V_low
+ 1.507010000e-07 V_low
+ 1.508000000e-07 V_low
+ 1.508010000e-07 V_low
+ 1.509000000e-07 V_low
+ 1.509010000e-07 V_hig
+ 1.510000000e-07 V_hig
+ 1.510010000e-07 V_hig
+ 1.511000000e-07 V_hig
+ 1.511010000e-07 V_hig
+ 1.512000000e-07 V_hig
+ 1.512010000e-07 V_hig
+ 1.513000000e-07 V_hig
+ 1.513010000e-07 V_hig
+ 1.514000000e-07 V_hig
+ 1.514010000e-07 V_hig
+ 1.515000000e-07 V_hig
+ 1.515010000e-07 V_hig
+ 1.516000000e-07 V_hig
+ 1.516010000e-07 V_hig
+ 1.517000000e-07 V_hig
+ 1.517010000e-07 V_hig
+ 1.518000000e-07 V_hig
+ 1.518010000e-07 V_hig
+ 1.519000000e-07 V_hig
+ 1.519010000e-07 V_low
+ 1.520000000e-07 V_low
+ 1.520010000e-07 V_low
+ 1.521000000e-07 V_low
+ 1.521010000e-07 V_low
+ 1.522000000e-07 V_low
+ 1.522010000e-07 V_low
+ 1.523000000e-07 V_low
+ 1.523010000e-07 V_low
+ 1.524000000e-07 V_low
+ 1.524010000e-07 V_low
+ 1.525000000e-07 V_low
+ 1.525010000e-07 V_low
+ 1.526000000e-07 V_low
+ 1.526010000e-07 V_low
+ 1.527000000e-07 V_low
+ 1.527010000e-07 V_low
+ 1.528000000e-07 V_low
+ 1.528010000e-07 V_low
+ 1.529000000e-07 V_low
+ 1.529010000e-07 V_hig
+ 1.530000000e-07 V_hig
+ 1.530010000e-07 V_hig
+ 1.531000000e-07 V_hig
+ 1.531010000e-07 V_hig
+ 1.532000000e-07 V_hig
+ 1.532010000e-07 V_hig
+ 1.533000000e-07 V_hig
+ 1.533010000e-07 V_hig
+ 1.534000000e-07 V_hig
+ 1.534010000e-07 V_hig
+ 1.535000000e-07 V_hig
+ 1.535010000e-07 V_hig
+ 1.536000000e-07 V_hig
+ 1.536010000e-07 V_hig
+ 1.537000000e-07 V_hig
+ 1.537010000e-07 V_hig
+ 1.538000000e-07 V_hig
+ 1.538010000e-07 V_hig
+ 1.539000000e-07 V_hig
+ 1.539010000e-07 V_low
+ 1.540000000e-07 V_low
+ 1.540010000e-07 V_low
+ 1.541000000e-07 V_low
+ 1.541010000e-07 V_low
+ 1.542000000e-07 V_low
+ 1.542010000e-07 V_low
+ 1.543000000e-07 V_low
+ 1.543010000e-07 V_low
+ 1.544000000e-07 V_low
+ 1.544010000e-07 V_low
+ 1.545000000e-07 V_low
+ 1.545010000e-07 V_low
+ 1.546000000e-07 V_low
+ 1.546010000e-07 V_low
+ 1.547000000e-07 V_low
+ 1.547010000e-07 V_low
+ 1.548000000e-07 V_low
+ 1.548010000e-07 V_low
+ 1.549000000e-07 V_low
+ 1.549010000e-07 V_low
+ 1.550000000e-07 V_low
+ 1.550010000e-07 V_low
+ 1.551000000e-07 V_low
+ 1.551010000e-07 V_low
+ 1.552000000e-07 V_low
+ 1.552010000e-07 V_low
+ 1.553000000e-07 V_low
+ 1.553010000e-07 V_low
+ 1.554000000e-07 V_low
+ 1.554010000e-07 V_low
+ 1.555000000e-07 V_low
+ 1.555010000e-07 V_low
+ 1.556000000e-07 V_low
+ 1.556010000e-07 V_low
+ 1.557000000e-07 V_low
+ 1.557010000e-07 V_low
+ 1.558000000e-07 V_low
+ 1.558010000e-07 V_low
+ 1.559000000e-07 V_low
+ 1.559010000e-07 V_hig
+ 1.560000000e-07 V_hig
+ 1.560010000e-07 V_hig
+ 1.561000000e-07 V_hig
+ 1.561010000e-07 V_hig
+ 1.562000000e-07 V_hig
+ 1.562010000e-07 V_hig
+ 1.563000000e-07 V_hig
+ 1.563010000e-07 V_hig
+ 1.564000000e-07 V_hig
+ 1.564010000e-07 V_hig
+ 1.565000000e-07 V_hig
+ 1.565010000e-07 V_hig
+ 1.566000000e-07 V_hig
+ 1.566010000e-07 V_hig
+ 1.567000000e-07 V_hig
+ 1.567010000e-07 V_hig
+ 1.568000000e-07 V_hig
+ 1.568010000e-07 V_hig
+ 1.569000000e-07 V_hig
+ 1.569010000e-07 V_hig
+ 1.570000000e-07 V_hig
+ 1.570010000e-07 V_hig
+ 1.571000000e-07 V_hig
+ 1.571010000e-07 V_hig
+ 1.572000000e-07 V_hig
+ 1.572010000e-07 V_hig
+ 1.573000000e-07 V_hig
+ 1.573010000e-07 V_hig
+ 1.574000000e-07 V_hig
+ 1.574010000e-07 V_hig
+ 1.575000000e-07 V_hig
+ 1.575010000e-07 V_hig
+ 1.576000000e-07 V_hig
+ 1.576010000e-07 V_hig
+ 1.577000000e-07 V_hig
+ 1.577010000e-07 V_hig
+ 1.578000000e-07 V_hig
+ 1.578010000e-07 V_hig
+ 1.579000000e-07 V_hig
+ 1.579010000e-07 V_hig
+ 1.580000000e-07 V_hig
+ 1.580010000e-07 V_hig
+ 1.581000000e-07 V_hig
+ 1.581010000e-07 V_hig
+ 1.582000000e-07 V_hig
+ 1.582010000e-07 V_hig
+ 1.583000000e-07 V_hig
+ 1.583010000e-07 V_hig
+ 1.584000000e-07 V_hig
+ 1.584010000e-07 V_hig
+ 1.585000000e-07 V_hig
+ 1.585010000e-07 V_hig
+ 1.586000000e-07 V_hig
+ 1.586010000e-07 V_hig
+ 1.587000000e-07 V_hig
+ 1.587010000e-07 V_hig
+ 1.588000000e-07 V_hig
+ 1.588010000e-07 V_hig
+ 1.589000000e-07 V_hig
+ 1.589010000e-07 V_hig
+ 1.590000000e-07 V_hig
+ 1.590010000e-07 V_hig
+ 1.591000000e-07 V_hig
+ 1.591010000e-07 V_hig
+ 1.592000000e-07 V_hig
+ 1.592010000e-07 V_hig
+ 1.593000000e-07 V_hig
+ 1.593010000e-07 V_hig
+ 1.594000000e-07 V_hig
+ 1.594010000e-07 V_hig
+ 1.595000000e-07 V_hig
+ 1.595010000e-07 V_hig
+ 1.596000000e-07 V_hig
+ 1.596010000e-07 V_hig
+ 1.597000000e-07 V_hig
+ 1.597010000e-07 V_hig
+ 1.598000000e-07 V_hig
+ 1.598010000e-07 V_hig
+ 1.599000000e-07 V_hig
+ 1.599010000e-07 V_hig
+ 1.600000000e-07 V_hig
+ 1.600010000e-07 V_hig
+ 1.601000000e-07 V_hig
+ 1.601010000e-07 V_hig
+ 1.602000000e-07 V_hig
+ 1.602010000e-07 V_hig
+ 1.603000000e-07 V_hig
+ 1.603010000e-07 V_hig
+ 1.604000000e-07 V_hig
+ 1.604010000e-07 V_hig
+ 1.605000000e-07 V_hig
+ 1.605010000e-07 V_hig
+ 1.606000000e-07 V_hig
+ 1.606010000e-07 V_hig
+ 1.607000000e-07 V_hig
+ 1.607010000e-07 V_hig
+ 1.608000000e-07 V_hig
+ 1.608010000e-07 V_hig
+ 1.609000000e-07 V_hig
+ 1.609010000e-07 V_low
+ 1.610000000e-07 V_low
+ 1.610010000e-07 V_low
+ 1.611000000e-07 V_low
+ 1.611010000e-07 V_low
+ 1.612000000e-07 V_low
+ 1.612010000e-07 V_low
+ 1.613000000e-07 V_low
+ 1.613010000e-07 V_low
+ 1.614000000e-07 V_low
+ 1.614010000e-07 V_low
+ 1.615000000e-07 V_low
+ 1.615010000e-07 V_low
+ 1.616000000e-07 V_low
+ 1.616010000e-07 V_low
+ 1.617000000e-07 V_low
+ 1.617010000e-07 V_low
+ 1.618000000e-07 V_low
+ 1.618010000e-07 V_low
+ 1.619000000e-07 V_low
+ 1.619010000e-07 V_low
+ 1.620000000e-07 V_low
+ 1.620010000e-07 V_low
+ 1.621000000e-07 V_low
+ 1.621010000e-07 V_low
+ 1.622000000e-07 V_low
+ 1.622010000e-07 V_low
+ 1.623000000e-07 V_low
+ 1.623010000e-07 V_low
+ 1.624000000e-07 V_low
+ 1.624010000e-07 V_low
+ 1.625000000e-07 V_low
+ 1.625010000e-07 V_low
+ 1.626000000e-07 V_low
+ 1.626010000e-07 V_low
+ 1.627000000e-07 V_low
+ 1.627010000e-07 V_low
+ 1.628000000e-07 V_low
+ 1.628010000e-07 V_low
+ 1.629000000e-07 V_low
+ 1.629010000e-07 V_hig
+ 1.630000000e-07 V_hig
+ 1.630010000e-07 V_hig
+ 1.631000000e-07 V_hig
+ 1.631010000e-07 V_hig
+ 1.632000000e-07 V_hig
+ 1.632010000e-07 V_hig
+ 1.633000000e-07 V_hig
+ 1.633010000e-07 V_hig
+ 1.634000000e-07 V_hig
+ 1.634010000e-07 V_hig
+ 1.635000000e-07 V_hig
+ 1.635010000e-07 V_hig
+ 1.636000000e-07 V_hig
+ 1.636010000e-07 V_hig
+ 1.637000000e-07 V_hig
+ 1.637010000e-07 V_hig
+ 1.638000000e-07 V_hig
+ 1.638010000e-07 V_hig
+ 1.639000000e-07 V_hig
+ 1.639010000e-07 V_hig
+ 1.640000000e-07 V_hig
+ 1.640010000e-07 V_hig
+ 1.641000000e-07 V_hig
+ 1.641010000e-07 V_hig
+ 1.642000000e-07 V_hig
+ 1.642010000e-07 V_hig
+ 1.643000000e-07 V_hig
+ 1.643010000e-07 V_hig
+ 1.644000000e-07 V_hig
+ 1.644010000e-07 V_hig
+ 1.645000000e-07 V_hig
+ 1.645010000e-07 V_hig
+ 1.646000000e-07 V_hig
+ 1.646010000e-07 V_hig
+ 1.647000000e-07 V_hig
+ 1.647010000e-07 V_hig
+ 1.648000000e-07 V_hig
+ 1.648010000e-07 V_hig
+ 1.649000000e-07 V_hig
+ 1.649010000e-07 V_hig
+ 1.650000000e-07 V_hig
+ 1.650010000e-07 V_hig
+ 1.651000000e-07 V_hig
+ 1.651010000e-07 V_hig
+ 1.652000000e-07 V_hig
+ 1.652010000e-07 V_hig
+ 1.653000000e-07 V_hig
+ 1.653010000e-07 V_hig
+ 1.654000000e-07 V_hig
+ 1.654010000e-07 V_hig
+ 1.655000000e-07 V_hig
+ 1.655010000e-07 V_hig
+ 1.656000000e-07 V_hig
+ 1.656010000e-07 V_hig
+ 1.657000000e-07 V_hig
+ 1.657010000e-07 V_hig
+ 1.658000000e-07 V_hig
+ 1.658010000e-07 V_hig
+ 1.659000000e-07 V_hig
+ 1.659010000e-07 V_hig
+ 1.660000000e-07 V_hig
+ 1.660010000e-07 V_hig
+ 1.661000000e-07 V_hig
+ 1.661010000e-07 V_hig
+ 1.662000000e-07 V_hig
+ 1.662010000e-07 V_hig
+ 1.663000000e-07 V_hig
+ 1.663010000e-07 V_hig
+ 1.664000000e-07 V_hig
+ 1.664010000e-07 V_hig
+ 1.665000000e-07 V_hig
+ 1.665010000e-07 V_hig
+ 1.666000000e-07 V_hig
+ 1.666010000e-07 V_hig
+ 1.667000000e-07 V_hig
+ 1.667010000e-07 V_hig
+ 1.668000000e-07 V_hig
+ 1.668010000e-07 V_hig
+ 1.669000000e-07 V_hig
+ 1.669010000e-07 V_hig
+ 1.670000000e-07 V_hig
+ 1.670010000e-07 V_hig
+ 1.671000000e-07 V_hig
+ 1.671010000e-07 V_hig
+ 1.672000000e-07 V_hig
+ 1.672010000e-07 V_hig
+ 1.673000000e-07 V_hig
+ 1.673010000e-07 V_hig
+ 1.674000000e-07 V_hig
+ 1.674010000e-07 V_hig
+ 1.675000000e-07 V_hig
+ 1.675010000e-07 V_hig
+ 1.676000000e-07 V_hig
+ 1.676010000e-07 V_hig
+ 1.677000000e-07 V_hig
+ 1.677010000e-07 V_hig
+ 1.678000000e-07 V_hig
+ 1.678010000e-07 V_hig
+ 1.679000000e-07 V_hig
+ 1.679010000e-07 V_low
+ 1.680000000e-07 V_low
+ 1.680010000e-07 V_low
+ 1.681000000e-07 V_low
+ 1.681010000e-07 V_low
+ 1.682000000e-07 V_low
+ 1.682010000e-07 V_low
+ 1.683000000e-07 V_low
+ 1.683010000e-07 V_low
+ 1.684000000e-07 V_low
+ 1.684010000e-07 V_low
+ 1.685000000e-07 V_low
+ 1.685010000e-07 V_low
+ 1.686000000e-07 V_low
+ 1.686010000e-07 V_low
+ 1.687000000e-07 V_low
+ 1.687010000e-07 V_low
+ 1.688000000e-07 V_low
+ 1.688010000e-07 V_low
+ 1.689000000e-07 V_low
+ 1.689010000e-07 V_low
+ 1.690000000e-07 V_low
+ 1.690010000e-07 V_low
+ 1.691000000e-07 V_low
+ 1.691010000e-07 V_low
+ 1.692000000e-07 V_low
+ 1.692010000e-07 V_low
+ 1.693000000e-07 V_low
+ 1.693010000e-07 V_low
+ 1.694000000e-07 V_low
+ 1.694010000e-07 V_low
+ 1.695000000e-07 V_low
+ 1.695010000e-07 V_low
+ 1.696000000e-07 V_low
+ 1.696010000e-07 V_low
+ 1.697000000e-07 V_low
+ 1.697010000e-07 V_low
+ 1.698000000e-07 V_low
+ 1.698010000e-07 V_low
+ 1.699000000e-07 V_low
+ 1.699010000e-07 V_hig
+ 1.700000000e-07 V_hig
+ 1.700010000e-07 V_hig
+ 1.701000000e-07 V_hig
+ 1.701010000e-07 V_hig
+ 1.702000000e-07 V_hig
+ 1.702010000e-07 V_hig
+ 1.703000000e-07 V_hig
+ 1.703010000e-07 V_hig
+ 1.704000000e-07 V_hig
+ 1.704010000e-07 V_hig
+ 1.705000000e-07 V_hig
+ 1.705010000e-07 V_hig
+ 1.706000000e-07 V_hig
+ 1.706010000e-07 V_hig
+ 1.707000000e-07 V_hig
+ 1.707010000e-07 V_hig
+ 1.708000000e-07 V_hig
+ 1.708010000e-07 V_hig
+ 1.709000000e-07 V_hig
+ 1.709010000e-07 V_low
+ 1.710000000e-07 V_low
+ 1.710010000e-07 V_low
+ 1.711000000e-07 V_low
+ 1.711010000e-07 V_low
+ 1.712000000e-07 V_low
+ 1.712010000e-07 V_low
+ 1.713000000e-07 V_low
+ 1.713010000e-07 V_low
+ 1.714000000e-07 V_low
+ 1.714010000e-07 V_low
+ 1.715000000e-07 V_low
+ 1.715010000e-07 V_low
+ 1.716000000e-07 V_low
+ 1.716010000e-07 V_low
+ 1.717000000e-07 V_low
+ 1.717010000e-07 V_low
+ 1.718000000e-07 V_low
+ 1.718010000e-07 V_low
+ 1.719000000e-07 V_low
+ 1.719010000e-07 V_hig
+ 1.720000000e-07 V_hig
+ 1.720010000e-07 V_hig
+ 1.721000000e-07 V_hig
+ 1.721010000e-07 V_hig
+ 1.722000000e-07 V_hig
+ 1.722010000e-07 V_hig
+ 1.723000000e-07 V_hig
+ 1.723010000e-07 V_hig
+ 1.724000000e-07 V_hig
+ 1.724010000e-07 V_hig
+ 1.725000000e-07 V_hig
+ 1.725010000e-07 V_hig
+ 1.726000000e-07 V_hig
+ 1.726010000e-07 V_hig
+ 1.727000000e-07 V_hig
+ 1.727010000e-07 V_hig
+ 1.728000000e-07 V_hig
+ 1.728010000e-07 V_hig
+ 1.729000000e-07 V_hig
+ 1.729010000e-07 V_hig
+ 1.730000000e-07 V_hig
+ 1.730010000e-07 V_hig
+ 1.731000000e-07 V_hig
+ 1.731010000e-07 V_hig
+ 1.732000000e-07 V_hig
+ 1.732010000e-07 V_hig
+ 1.733000000e-07 V_hig
+ 1.733010000e-07 V_hig
+ 1.734000000e-07 V_hig
+ 1.734010000e-07 V_hig
+ 1.735000000e-07 V_hig
+ 1.735010000e-07 V_hig
+ 1.736000000e-07 V_hig
+ 1.736010000e-07 V_hig
+ 1.737000000e-07 V_hig
+ 1.737010000e-07 V_hig
+ 1.738000000e-07 V_hig
+ 1.738010000e-07 V_hig
+ 1.739000000e-07 V_hig
+ 1.739010000e-07 V_low
+ 1.740000000e-07 V_low
+ 1.740010000e-07 V_low
+ 1.741000000e-07 V_low
+ 1.741010000e-07 V_low
+ 1.742000000e-07 V_low
+ 1.742010000e-07 V_low
+ 1.743000000e-07 V_low
+ 1.743010000e-07 V_low
+ 1.744000000e-07 V_low
+ 1.744010000e-07 V_low
+ 1.745000000e-07 V_low
+ 1.745010000e-07 V_low
+ 1.746000000e-07 V_low
+ 1.746010000e-07 V_low
+ 1.747000000e-07 V_low
+ 1.747010000e-07 V_low
+ 1.748000000e-07 V_low
+ 1.748010000e-07 V_low
+ 1.749000000e-07 V_low
+ 1.749010000e-07 V_low
+ 1.750000000e-07 V_low
+ 1.750010000e-07 V_low
+ 1.751000000e-07 V_low
+ 1.751010000e-07 V_low
+ 1.752000000e-07 V_low
+ 1.752010000e-07 V_low
+ 1.753000000e-07 V_low
+ 1.753010000e-07 V_low
+ 1.754000000e-07 V_low
+ 1.754010000e-07 V_low
+ 1.755000000e-07 V_low
+ 1.755010000e-07 V_low
+ 1.756000000e-07 V_low
+ 1.756010000e-07 V_low
+ 1.757000000e-07 V_low
+ 1.757010000e-07 V_low
+ 1.758000000e-07 V_low
+ 1.758010000e-07 V_low
+ 1.759000000e-07 V_low
+ 1.759010000e-07 V_low
+ 1.760000000e-07 V_low
+ 1.760010000e-07 V_low
+ 1.761000000e-07 V_low
+ 1.761010000e-07 V_low
+ 1.762000000e-07 V_low
+ 1.762010000e-07 V_low
+ 1.763000000e-07 V_low
+ 1.763010000e-07 V_low
+ 1.764000000e-07 V_low
+ 1.764010000e-07 V_low
+ 1.765000000e-07 V_low
+ 1.765010000e-07 V_low
+ 1.766000000e-07 V_low
+ 1.766010000e-07 V_low
+ 1.767000000e-07 V_low
+ 1.767010000e-07 V_low
+ 1.768000000e-07 V_low
+ 1.768010000e-07 V_low
+ 1.769000000e-07 V_low
+ 1.769010000e-07 V_hig
+ 1.770000000e-07 V_hig
+ 1.770010000e-07 V_hig
+ 1.771000000e-07 V_hig
+ 1.771010000e-07 V_hig
+ 1.772000000e-07 V_hig
+ 1.772010000e-07 V_hig
+ 1.773000000e-07 V_hig
+ 1.773010000e-07 V_hig
+ 1.774000000e-07 V_hig
+ 1.774010000e-07 V_hig
+ 1.775000000e-07 V_hig
+ 1.775010000e-07 V_hig
+ 1.776000000e-07 V_hig
+ 1.776010000e-07 V_hig
+ 1.777000000e-07 V_hig
+ 1.777010000e-07 V_hig
+ 1.778000000e-07 V_hig
+ 1.778010000e-07 V_hig
+ 1.779000000e-07 V_hig
+ 1.779010000e-07 V_low
+ 1.780000000e-07 V_low
+ 1.780010000e-07 V_low
+ 1.781000000e-07 V_low
+ 1.781010000e-07 V_low
+ 1.782000000e-07 V_low
+ 1.782010000e-07 V_low
+ 1.783000000e-07 V_low
+ 1.783010000e-07 V_low
+ 1.784000000e-07 V_low
+ 1.784010000e-07 V_low
+ 1.785000000e-07 V_low
+ 1.785010000e-07 V_low
+ 1.786000000e-07 V_low
+ 1.786010000e-07 V_low
+ 1.787000000e-07 V_low
+ 1.787010000e-07 V_low
+ 1.788000000e-07 V_low
+ 1.788010000e-07 V_low
+ 1.789000000e-07 V_low
+ 1.789010000e-07 V_hig
+ 1.790000000e-07 V_hig
+ 1.790010000e-07 V_hig
+ 1.791000000e-07 V_hig
+ 1.791010000e-07 V_hig
+ 1.792000000e-07 V_hig
+ 1.792010000e-07 V_hig
+ 1.793000000e-07 V_hig
+ 1.793010000e-07 V_hig
+ 1.794000000e-07 V_hig
+ 1.794010000e-07 V_hig
+ 1.795000000e-07 V_hig
+ 1.795010000e-07 V_hig
+ 1.796000000e-07 V_hig
+ 1.796010000e-07 V_hig
+ 1.797000000e-07 V_hig
+ 1.797010000e-07 V_hig
+ 1.798000000e-07 V_hig
+ 1.798010000e-07 V_hig
+ 1.799000000e-07 V_hig
+ 1.799010000e-07 V_low
+ 1.800000000e-07 V_low
+ 1.800010000e-07 V_low
+ 1.801000000e-07 V_low
+ 1.801010000e-07 V_low
+ 1.802000000e-07 V_low
+ 1.802010000e-07 V_low
+ 1.803000000e-07 V_low
+ 1.803010000e-07 V_low
+ 1.804000000e-07 V_low
+ 1.804010000e-07 V_low
+ 1.805000000e-07 V_low
+ 1.805010000e-07 V_low
+ 1.806000000e-07 V_low
+ 1.806010000e-07 V_low
+ 1.807000000e-07 V_low
+ 1.807010000e-07 V_low
+ 1.808000000e-07 V_low
+ 1.808010000e-07 V_low
+ 1.809000000e-07 V_low
+ 1.809010000e-07 V_low
+ 1.810000000e-07 V_low
+ 1.810010000e-07 V_low
+ 1.811000000e-07 V_low
+ 1.811010000e-07 V_low
+ 1.812000000e-07 V_low
+ 1.812010000e-07 V_low
+ 1.813000000e-07 V_low
+ 1.813010000e-07 V_low
+ 1.814000000e-07 V_low
+ 1.814010000e-07 V_low
+ 1.815000000e-07 V_low
+ 1.815010000e-07 V_low
+ 1.816000000e-07 V_low
+ 1.816010000e-07 V_low
+ 1.817000000e-07 V_low
+ 1.817010000e-07 V_low
+ 1.818000000e-07 V_low
+ 1.818010000e-07 V_low
+ 1.819000000e-07 V_low
+ 1.819010000e-07 V_low
+ 1.820000000e-07 V_low
+ 1.820010000e-07 V_low
+ 1.821000000e-07 V_low
+ 1.821010000e-07 V_low
+ 1.822000000e-07 V_low
+ 1.822010000e-07 V_low
+ 1.823000000e-07 V_low
+ 1.823010000e-07 V_low
+ 1.824000000e-07 V_low
+ 1.824010000e-07 V_low
+ 1.825000000e-07 V_low
+ 1.825010000e-07 V_low
+ 1.826000000e-07 V_low
+ 1.826010000e-07 V_low
+ 1.827000000e-07 V_low
+ 1.827010000e-07 V_low
+ 1.828000000e-07 V_low
+ 1.828010000e-07 V_low
+ 1.829000000e-07 V_low
+ 1.829010000e-07 V_hig
+ 1.830000000e-07 V_hig
+ 1.830010000e-07 V_hig
+ 1.831000000e-07 V_hig
+ 1.831010000e-07 V_hig
+ 1.832000000e-07 V_hig
+ 1.832010000e-07 V_hig
+ 1.833000000e-07 V_hig
+ 1.833010000e-07 V_hig
+ 1.834000000e-07 V_hig
+ 1.834010000e-07 V_hig
+ 1.835000000e-07 V_hig
+ 1.835010000e-07 V_hig
+ 1.836000000e-07 V_hig
+ 1.836010000e-07 V_hig
+ 1.837000000e-07 V_hig
+ 1.837010000e-07 V_hig
+ 1.838000000e-07 V_hig
+ 1.838010000e-07 V_hig
+ 1.839000000e-07 V_hig
+ 1.839010000e-07 V_hig
+ 1.840000000e-07 V_hig
+ 1.840010000e-07 V_hig
+ 1.841000000e-07 V_hig
+ 1.841010000e-07 V_hig
+ 1.842000000e-07 V_hig
+ 1.842010000e-07 V_hig
+ 1.843000000e-07 V_hig
+ 1.843010000e-07 V_hig
+ 1.844000000e-07 V_hig
+ 1.844010000e-07 V_hig
+ 1.845000000e-07 V_hig
+ 1.845010000e-07 V_hig
+ 1.846000000e-07 V_hig
+ 1.846010000e-07 V_hig
+ 1.847000000e-07 V_hig
+ 1.847010000e-07 V_hig
+ 1.848000000e-07 V_hig
+ 1.848010000e-07 V_hig
+ 1.849000000e-07 V_hig
+ 1.849010000e-07 V_low
+ 1.850000000e-07 V_low
+ 1.850010000e-07 V_low
+ 1.851000000e-07 V_low
+ 1.851010000e-07 V_low
+ 1.852000000e-07 V_low
+ 1.852010000e-07 V_low
+ 1.853000000e-07 V_low
+ 1.853010000e-07 V_low
+ 1.854000000e-07 V_low
+ 1.854010000e-07 V_low
+ 1.855000000e-07 V_low
+ 1.855010000e-07 V_low
+ 1.856000000e-07 V_low
+ 1.856010000e-07 V_low
+ 1.857000000e-07 V_low
+ 1.857010000e-07 V_low
+ 1.858000000e-07 V_low
+ 1.858010000e-07 V_low
+ 1.859000000e-07 V_low
+ 1.859010000e-07 V_low
+ 1.860000000e-07 V_low
+ 1.860010000e-07 V_low
+ 1.861000000e-07 V_low
+ 1.861010000e-07 V_low
+ 1.862000000e-07 V_low
+ 1.862010000e-07 V_low
+ 1.863000000e-07 V_low
+ 1.863010000e-07 V_low
+ 1.864000000e-07 V_low
+ 1.864010000e-07 V_low
+ 1.865000000e-07 V_low
+ 1.865010000e-07 V_low
+ 1.866000000e-07 V_low
+ 1.866010000e-07 V_low
+ 1.867000000e-07 V_low
+ 1.867010000e-07 V_low
+ 1.868000000e-07 V_low
+ 1.868010000e-07 V_low
+ 1.869000000e-07 V_low
+ 1.869010000e-07 V_low
+ 1.870000000e-07 V_low
+ 1.870010000e-07 V_low
+ 1.871000000e-07 V_low
+ 1.871010000e-07 V_low
+ 1.872000000e-07 V_low
+ 1.872010000e-07 V_low
+ 1.873000000e-07 V_low
+ 1.873010000e-07 V_low
+ 1.874000000e-07 V_low
+ 1.874010000e-07 V_low
+ 1.875000000e-07 V_low
+ 1.875010000e-07 V_low
+ 1.876000000e-07 V_low
+ 1.876010000e-07 V_low
+ 1.877000000e-07 V_low
+ 1.877010000e-07 V_low
+ 1.878000000e-07 V_low
+ 1.878010000e-07 V_low
+ 1.879000000e-07 V_low
+ 1.879010000e-07 V_low
+ 1.880000000e-07 V_low
+ 1.880010000e-07 V_low
+ 1.881000000e-07 V_low
+ 1.881010000e-07 V_low
+ 1.882000000e-07 V_low
+ 1.882010000e-07 V_low
+ 1.883000000e-07 V_low
+ 1.883010000e-07 V_low
+ 1.884000000e-07 V_low
+ 1.884010000e-07 V_low
+ 1.885000000e-07 V_low
+ 1.885010000e-07 V_low
+ 1.886000000e-07 V_low
+ 1.886010000e-07 V_low
+ 1.887000000e-07 V_low
+ 1.887010000e-07 V_low
+ 1.888000000e-07 V_low
+ 1.888010000e-07 V_low
+ 1.889000000e-07 V_low
+ 1.889010000e-07 V_hig
+ 1.890000000e-07 V_hig
+ 1.890010000e-07 V_hig
+ 1.891000000e-07 V_hig
+ 1.891010000e-07 V_hig
+ 1.892000000e-07 V_hig
+ 1.892010000e-07 V_hig
+ 1.893000000e-07 V_hig
+ 1.893010000e-07 V_hig
+ 1.894000000e-07 V_hig
+ 1.894010000e-07 V_hig
+ 1.895000000e-07 V_hig
+ 1.895010000e-07 V_hig
+ 1.896000000e-07 V_hig
+ 1.896010000e-07 V_hig
+ 1.897000000e-07 V_hig
+ 1.897010000e-07 V_hig
+ 1.898000000e-07 V_hig
+ 1.898010000e-07 V_hig
+ 1.899000000e-07 V_hig
+ 1.899010000e-07 V_hig
+ 1.900000000e-07 V_hig
+ 1.900010000e-07 V_hig
+ 1.901000000e-07 V_hig
+ 1.901010000e-07 V_hig
+ 1.902000000e-07 V_hig
+ 1.902010000e-07 V_hig
+ 1.903000000e-07 V_hig
+ 1.903010000e-07 V_hig
+ 1.904000000e-07 V_hig
+ 1.904010000e-07 V_hig
+ 1.905000000e-07 V_hig
+ 1.905010000e-07 V_hig
+ 1.906000000e-07 V_hig
+ 1.906010000e-07 V_hig
+ 1.907000000e-07 V_hig
+ 1.907010000e-07 V_hig
+ 1.908000000e-07 V_hig
+ 1.908010000e-07 V_hig
+ 1.909000000e-07 V_hig
+ 1.909010000e-07 V_low
+ 1.910000000e-07 V_low
+ 1.910010000e-07 V_low
+ 1.911000000e-07 V_low
+ 1.911010000e-07 V_low
+ 1.912000000e-07 V_low
+ 1.912010000e-07 V_low
+ 1.913000000e-07 V_low
+ 1.913010000e-07 V_low
+ 1.914000000e-07 V_low
+ 1.914010000e-07 V_low
+ 1.915000000e-07 V_low
+ 1.915010000e-07 V_low
+ 1.916000000e-07 V_low
+ 1.916010000e-07 V_low
+ 1.917000000e-07 V_low
+ 1.917010000e-07 V_low
+ 1.918000000e-07 V_low
+ 1.918010000e-07 V_low
+ 1.919000000e-07 V_low
+ 1.919010000e-07 V_low
+ 1.920000000e-07 V_low
+ 1.920010000e-07 V_low
+ 1.921000000e-07 V_low
+ 1.921010000e-07 V_low
+ 1.922000000e-07 V_low
+ 1.922010000e-07 V_low
+ 1.923000000e-07 V_low
+ 1.923010000e-07 V_low
+ 1.924000000e-07 V_low
+ 1.924010000e-07 V_low
+ 1.925000000e-07 V_low
+ 1.925010000e-07 V_low
+ 1.926000000e-07 V_low
+ 1.926010000e-07 V_low
+ 1.927000000e-07 V_low
+ 1.927010000e-07 V_low
+ 1.928000000e-07 V_low
+ 1.928010000e-07 V_low
+ 1.929000000e-07 V_low
+ 1.929010000e-07 V_low
+ 1.930000000e-07 V_low
+ 1.930010000e-07 V_low
+ 1.931000000e-07 V_low
+ 1.931010000e-07 V_low
+ 1.932000000e-07 V_low
+ 1.932010000e-07 V_low
+ 1.933000000e-07 V_low
+ 1.933010000e-07 V_low
+ 1.934000000e-07 V_low
+ 1.934010000e-07 V_low
+ 1.935000000e-07 V_low
+ 1.935010000e-07 V_low
+ 1.936000000e-07 V_low
+ 1.936010000e-07 V_low
+ 1.937000000e-07 V_low
+ 1.937010000e-07 V_low
+ 1.938000000e-07 V_low
+ 1.938010000e-07 V_low
+ 1.939000000e-07 V_low
+ 1.939010000e-07 V_hig
+ 1.940000000e-07 V_hig
+ 1.940010000e-07 V_hig
+ 1.941000000e-07 V_hig
+ 1.941010000e-07 V_hig
+ 1.942000000e-07 V_hig
+ 1.942010000e-07 V_hig
+ 1.943000000e-07 V_hig
+ 1.943010000e-07 V_hig
+ 1.944000000e-07 V_hig
+ 1.944010000e-07 V_hig
+ 1.945000000e-07 V_hig
+ 1.945010000e-07 V_hig
+ 1.946000000e-07 V_hig
+ 1.946010000e-07 V_hig
+ 1.947000000e-07 V_hig
+ 1.947010000e-07 V_hig
+ 1.948000000e-07 V_hig
+ 1.948010000e-07 V_hig
+ 1.949000000e-07 V_hig
+ 1.949010000e-07 V_hig
+ 1.950000000e-07 V_hig
+ 1.950010000e-07 V_hig
+ 1.951000000e-07 V_hig
+ 1.951010000e-07 V_hig
+ 1.952000000e-07 V_hig
+ 1.952010000e-07 V_hig
+ 1.953000000e-07 V_hig
+ 1.953010000e-07 V_hig
+ 1.954000000e-07 V_hig
+ 1.954010000e-07 V_hig
+ 1.955000000e-07 V_hig
+ 1.955010000e-07 V_hig
+ 1.956000000e-07 V_hig
+ 1.956010000e-07 V_hig
+ 1.957000000e-07 V_hig
+ 1.957010000e-07 V_hig
+ 1.958000000e-07 V_hig
+ 1.958010000e-07 V_hig
+ 1.959000000e-07 V_hig
+ 1.959010000e-07 V_low
+ 1.960000000e-07 V_low
+ 1.960010000e-07 V_low
+ 1.961000000e-07 V_low
+ 1.961010000e-07 V_low
+ 1.962000000e-07 V_low
+ 1.962010000e-07 V_low
+ 1.963000000e-07 V_low
+ 1.963010000e-07 V_low
+ 1.964000000e-07 V_low
+ 1.964010000e-07 V_low
+ 1.965000000e-07 V_low
+ 1.965010000e-07 V_low
+ 1.966000000e-07 V_low
+ 1.966010000e-07 V_low
+ 1.967000000e-07 V_low
+ 1.967010000e-07 V_low
+ 1.968000000e-07 V_low
+ 1.968010000e-07 V_low
+ 1.969000000e-07 V_low
+ 1.969010000e-07 V_hig
+ 1.970000000e-07 V_hig
+ 1.970010000e-07 V_hig
+ 1.971000000e-07 V_hig
+ 1.971010000e-07 V_hig
+ 1.972000000e-07 V_hig
+ 1.972010000e-07 V_hig
+ 1.973000000e-07 V_hig
+ 1.973010000e-07 V_hig
+ 1.974000000e-07 V_hig
+ 1.974010000e-07 V_hig
+ 1.975000000e-07 V_hig
+ 1.975010000e-07 V_hig
+ 1.976000000e-07 V_hig
+ 1.976010000e-07 V_hig
+ 1.977000000e-07 V_hig
+ 1.977010000e-07 V_hig
+ 1.978000000e-07 V_hig
+ 1.978010000e-07 V_hig
+ 1.979000000e-07 V_hig
+ 1.979010000e-07 V_hig
+ 1.980000000e-07 V_hig
+ 1.980010000e-07 V_hig
+ 1.981000000e-07 V_hig
+ 1.981010000e-07 V_hig
+ 1.982000000e-07 V_hig
+ 1.982010000e-07 V_hig
+ 1.983000000e-07 V_hig
+ 1.983010000e-07 V_hig
+ 1.984000000e-07 V_hig
+ 1.984010000e-07 V_hig
+ 1.985000000e-07 V_hig
+ 1.985010000e-07 V_hig
+ 1.986000000e-07 V_hig
+ 1.986010000e-07 V_hig
+ 1.987000000e-07 V_hig
+ 1.987010000e-07 V_hig
+ 1.988000000e-07 V_hig
+ 1.988010000e-07 V_hig
+ 1.989000000e-07 V_hig
+ 1.989010000e-07 V_low
+ 1.990000000e-07 V_low
+ 1.990010000e-07 V_low
+ 1.991000000e-07 V_low
+ 1.991010000e-07 V_low
+ 1.992000000e-07 V_low
+ 1.992010000e-07 V_low
+ 1.993000000e-07 V_low
+ 1.993010000e-07 V_low
+ 1.994000000e-07 V_low
+ 1.994010000e-07 V_low
+ 1.995000000e-07 V_low
+ 1.995010000e-07 V_low
+ 1.996000000e-07 V_low
+ 1.996010000e-07 V_low
+ 1.997000000e-07 V_low
+ 1.997010000e-07 V_low
+ 1.998000000e-07 V_low
+ 1.998010000e-07 V_low
+ 1.999000000e-07 V_low
+ 1.999010000e-07 V_low
+ 2.000000000e-07 V_low
+ 2.000010000e-07 V_low
+ 2.001000000e-07 V_low
+ 2.001010000e-07 V_low
+ 2.002000000e-07 V_low
+ 2.002010000e-07 V_low
+ 2.003000000e-07 V_low
+ 2.003010000e-07 V_low
+ 2.004000000e-07 V_low
+ 2.004010000e-07 V_low
+ 2.005000000e-07 V_low
+ 2.005010000e-07 V_low
+ 2.006000000e-07 V_low
+ 2.006010000e-07 V_low
+ 2.007000000e-07 V_low
+ 2.007010000e-07 V_low
+ 2.008000000e-07 V_low
+ 2.008010000e-07 V_low
+ 2.009000000e-07 V_low
+ 2.009010000e-07 V_low
+ 2.010000000e-07 V_low
+ 2.010010000e-07 V_low
+ 2.011000000e-07 V_low
+ 2.011010000e-07 V_low
+ 2.012000000e-07 V_low
+ 2.012010000e-07 V_low
+ 2.013000000e-07 V_low
+ 2.013010000e-07 V_low
+ 2.014000000e-07 V_low
+ 2.014010000e-07 V_low
+ 2.015000000e-07 V_low
+ 2.015010000e-07 V_low
+ 2.016000000e-07 V_low
+ 2.016010000e-07 V_low
+ 2.017000000e-07 V_low
+ 2.017010000e-07 V_low
+ 2.018000000e-07 V_low
+ 2.018010000e-07 V_low
+ 2.019000000e-07 V_low
+ 2.019010000e-07 V_low
+ 2.020000000e-07 V_low
+ 2.020010000e-07 V_low
+ 2.021000000e-07 V_low
+ 2.021010000e-07 V_low
+ 2.022000000e-07 V_low
+ 2.022010000e-07 V_low
+ 2.023000000e-07 V_low
+ 2.023010000e-07 V_low
+ 2.024000000e-07 V_low
+ 2.024010000e-07 V_low
+ 2.025000000e-07 V_low
+ 2.025010000e-07 V_low
+ 2.026000000e-07 V_low
+ 2.026010000e-07 V_low
+ 2.027000000e-07 V_low
+ 2.027010000e-07 V_low
+ 2.028000000e-07 V_low
+ 2.028010000e-07 V_low
+ 2.029000000e-07 V_low
+ 2.029010000e-07 V_low
+ 2.030000000e-07 V_low
+ 2.030010000e-07 V_low
+ 2.031000000e-07 V_low
+ 2.031010000e-07 V_low
+ 2.032000000e-07 V_low
+ 2.032010000e-07 V_low
+ 2.033000000e-07 V_low
+ 2.033010000e-07 V_low
+ 2.034000000e-07 V_low
+ 2.034010000e-07 V_low
+ 2.035000000e-07 V_low
+ 2.035010000e-07 V_low
+ 2.036000000e-07 V_low
+ 2.036010000e-07 V_low
+ 2.037000000e-07 V_low
+ 2.037010000e-07 V_low
+ 2.038000000e-07 V_low
+ 2.038010000e-07 V_low
+ 2.039000000e-07 V_low
+ 2.039010000e-07 V_hig
+ 2.040000000e-07 V_hig
+ 2.040010000e-07 V_hig
+ 2.041000000e-07 V_hig
+ 2.041010000e-07 V_hig
+ 2.042000000e-07 V_hig
+ 2.042010000e-07 V_hig
+ 2.043000000e-07 V_hig
+ 2.043010000e-07 V_hig
+ 2.044000000e-07 V_hig
+ 2.044010000e-07 V_hig
+ 2.045000000e-07 V_hig
+ 2.045010000e-07 V_hig
+ 2.046000000e-07 V_hig
+ 2.046010000e-07 V_hig
+ 2.047000000e-07 V_hig
+ 2.047010000e-07 V_hig
+ 2.048000000e-07 V_hig
+ 2.048010000e-07 V_hig
+ 2.049000000e-07 V_hig
+ 2.049010000e-07 V_hig
+ 2.050000000e-07 V_hig
+ 2.050010000e-07 V_hig
+ 2.051000000e-07 V_hig
+ 2.051010000e-07 V_hig
+ 2.052000000e-07 V_hig
+ 2.052010000e-07 V_hig
+ 2.053000000e-07 V_hig
+ 2.053010000e-07 V_hig
+ 2.054000000e-07 V_hig
+ 2.054010000e-07 V_hig
+ 2.055000000e-07 V_hig
+ 2.055010000e-07 V_hig
+ 2.056000000e-07 V_hig
+ 2.056010000e-07 V_hig
+ 2.057000000e-07 V_hig
+ 2.057010000e-07 V_hig
+ 2.058000000e-07 V_hig
+ 2.058010000e-07 V_hig
+ 2.059000000e-07 V_hig
+ 2.059010000e-07 V_low
+ 2.060000000e-07 V_low
+ 2.060010000e-07 V_low
+ 2.061000000e-07 V_low
+ 2.061010000e-07 V_low
+ 2.062000000e-07 V_low
+ 2.062010000e-07 V_low
+ 2.063000000e-07 V_low
+ 2.063010000e-07 V_low
+ 2.064000000e-07 V_low
+ 2.064010000e-07 V_low
+ 2.065000000e-07 V_low
+ 2.065010000e-07 V_low
+ 2.066000000e-07 V_low
+ 2.066010000e-07 V_low
+ 2.067000000e-07 V_low
+ 2.067010000e-07 V_low
+ 2.068000000e-07 V_low
+ 2.068010000e-07 V_low
+ 2.069000000e-07 V_low
+ 2.069010000e-07 V_hig
+ 2.070000000e-07 V_hig
+ 2.070010000e-07 V_hig
+ 2.071000000e-07 V_hig
+ 2.071010000e-07 V_hig
+ 2.072000000e-07 V_hig
+ 2.072010000e-07 V_hig
+ 2.073000000e-07 V_hig
+ 2.073010000e-07 V_hig
+ 2.074000000e-07 V_hig
+ 2.074010000e-07 V_hig
+ 2.075000000e-07 V_hig
+ 2.075010000e-07 V_hig
+ 2.076000000e-07 V_hig
+ 2.076010000e-07 V_hig
+ 2.077000000e-07 V_hig
+ 2.077010000e-07 V_hig
+ 2.078000000e-07 V_hig
+ 2.078010000e-07 V_hig
+ 2.079000000e-07 V_hig
+ 2.079010000e-07 V_hig
+ 2.080000000e-07 V_hig
+ 2.080010000e-07 V_hig
+ 2.081000000e-07 V_hig
+ 2.081010000e-07 V_hig
+ 2.082000000e-07 V_hig
+ 2.082010000e-07 V_hig
+ 2.083000000e-07 V_hig
+ 2.083010000e-07 V_hig
+ 2.084000000e-07 V_hig
+ 2.084010000e-07 V_hig
+ 2.085000000e-07 V_hig
+ 2.085010000e-07 V_hig
+ 2.086000000e-07 V_hig
+ 2.086010000e-07 V_hig
+ 2.087000000e-07 V_hig
+ 2.087010000e-07 V_hig
+ 2.088000000e-07 V_hig
+ 2.088010000e-07 V_hig
+ 2.089000000e-07 V_hig
+ 2.089010000e-07 V_hig
+ 2.090000000e-07 V_hig
+ 2.090010000e-07 V_hig
+ 2.091000000e-07 V_hig
+ 2.091010000e-07 V_hig
+ 2.092000000e-07 V_hig
+ 2.092010000e-07 V_hig
+ 2.093000000e-07 V_hig
+ 2.093010000e-07 V_hig
+ 2.094000000e-07 V_hig
+ 2.094010000e-07 V_hig
+ 2.095000000e-07 V_hig
+ 2.095010000e-07 V_hig
+ 2.096000000e-07 V_hig
+ 2.096010000e-07 V_hig
+ 2.097000000e-07 V_hig
+ 2.097010000e-07 V_hig
+ 2.098000000e-07 V_hig
+ 2.098010000e-07 V_hig
+ 2.099000000e-07 V_hig
+ 2.099010000e-07 V_hig
+ 2.100000000e-07 V_hig
+ 2.100010000e-07 V_hig
+ 2.101000000e-07 V_hig
+ 2.101010000e-07 V_hig
+ 2.102000000e-07 V_hig
+ 2.102010000e-07 V_hig
+ 2.103000000e-07 V_hig
+ 2.103010000e-07 V_hig
+ 2.104000000e-07 V_hig
+ 2.104010000e-07 V_hig
+ 2.105000000e-07 V_hig
+ 2.105010000e-07 V_hig
+ 2.106000000e-07 V_hig
+ 2.106010000e-07 V_hig
+ 2.107000000e-07 V_hig
+ 2.107010000e-07 V_hig
+ 2.108000000e-07 V_hig
+ 2.108010000e-07 V_hig
+ 2.109000000e-07 V_hig
+ 2.109010000e-07 V_low
+ 2.110000000e-07 V_low
+ 2.110010000e-07 V_low
+ 2.111000000e-07 V_low
+ 2.111010000e-07 V_low
+ 2.112000000e-07 V_low
+ 2.112010000e-07 V_low
+ 2.113000000e-07 V_low
+ 2.113010000e-07 V_low
+ 2.114000000e-07 V_low
+ 2.114010000e-07 V_low
+ 2.115000000e-07 V_low
+ 2.115010000e-07 V_low
+ 2.116000000e-07 V_low
+ 2.116010000e-07 V_low
+ 2.117000000e-07 V_low
+ 2.117010000e-07 V_low
+ 2.118000000e-07 V_low
+ 2.118010000e-07 V_low
+ 2.119000000e-07 V_low
+ 2.119010000e-07 V_low
+ 2.120000000e-07 V_low
+ 2.120010000e-07 V_low
+ 2.121000000e-07 V_low
+ 2.121010000e-07 V_low
+ 2.122000000e-07 V_low
+ 2.122010000e-07 V_low
+ 2.123000000e-07 V_low
+ 2.123010000e-07 V_low
+ 2.124000000e-07 V_low
+ 2.124010000e-07 V_low
+ 2.125000000e-07 V_low
+ 2.125010000e-07 V_low
+ 2.126000000e-07 V_low
+ 2.126010000e-07 V_low
+ 2.127000000e-07 V_low
+ 2.127010000e-07 V_low
+ 2.128000000e-07 V_low
+ 2.128010000e-07 V_low
+ 2.129000000e-07 V_low
+ 2.129010000e-07 V_hig
+ 2.130000000e-07 V_hig
+ 2.130010000e-07 V_hig
+ 2.131000000e-07 V_hig
+ 2.131010000e-07 V_hig
+ 2.132000000e-07 V_hig
+ 2.132010000e-07 V_hig
+ 2.133000000e-07 V_hig
+ 2.133010000e-07 V_hig
+ 2.134000000e-07 V_hig
+ 2.134010000e-07 V_hig
+ 2.135000000e-07 V_hig
+ 2.135010000e-07 V_hig
+ 2.136000000e-07 V_hig
+ 2.136010000e-07 V_hig
+ 2.137000000e-07 V_hig
+ 2.137010000e-07 V_hig
+ 2.138000000e-07 V_hig
+ 2.138010000e-07 V_hig
+ 2.139000000e-07 V_hig
+ 2.139010000e-07 V_hig
+ 2.140000000e-07 V_hig
+ 2.140010000e-07 V_hig
+ 2.141000000e-07 V_hig
+ 2.141010000e-07 V_hig
+ 2.142000000e-07 V_hig
+ 2.142010000e-07 V_hig
+ 2.143000000e-07 V_hig
+ 2.143010000e-07 V_hig
+ 2.144000000e-07 V_hig
+ 2.144010000e-07 V_hig
+ 2.145000000e-07 V_hig
+ 2.145010000e-07 V_hig
+ 2.146000000e-07 V_hig
+ 2.146010000e-07 V_hig
+ 2.147000000e-07 V_hig
+ 2.147010000e-07 V_hig
+ 2.148000000e-07 V_hig
+ 2.148010000e-07 V_hig
+ 2.149000000e-07 V_hig
+ 2.149010000e-07 V_low
+ 2.150000000e-07 V_low
+ 2.150010000e-07 V_low
+ 2.151000000e-07 V_low
+ 2.151010000e-07 V_low
+ 2.152000000e-07 V_low
+ 2.152010000e-07 V_low
+ 2.153000000e-07 V_low
+ 2.153010000e-07 V_low
+ 2.154000000e-07 V_low
+ 2.154010000e-07 V_low
+ 2.155000000e-07 V_low
+ 2.155010000e-07 V_low
+ 2.156000000e-07 V_low
+ 2.156010000e-07 V_low
+ 2.157000000e-07 V_low
+ 2.157010000e-07 V_low
+ 2.158000000e-07 V_low
+ 2.158010000e-07 V_low
+ 2.159000000e-07 V_low
+ 2.159010000e-07 V_hig
+ 2.160000000e-07 V_hig
+ 2.160010000e-07 V_hig
+ 2.161000000e-07 V_hig
+ 2.161010000e-07 V_hig
+ 2.162000000e-07 V_hig
+ 2.162010000e-07 V_hig
+ 2.163000000e-07 V_hig
+ 2.163010000e-07 V_hig
+ 2.164000000e-07 V_hig
+ 2.164010000e-07 V_hig
+ 2.165000000e-07 V_hig
+ 2.165010000e-07 V_hig
+ 2.166000000e-07 V_hig
+ 2.166010000e-07 V_hig
+ 2.167000000e-07 V_hig
+ 2.167010000e-07 V_hig
+ 2.168000000e-07 V_hig
+ 2.168010000e-07 V_hig
+ 2.169000000e-07 V_hig
+ 2.169010000e-07 V_hig
+ 2.170000000e-07 V_hig
+ 2.170010000e-07 V_hig
+ 2.171000000e-07 V_hig
+ 2.171010000e-07 V_hig
+ 2.172000000e-07 V_hig
+ 2.172010000e-07 V_hig
+ 2.173000000e-07 V_hig
+ 2.173010000e-07 V_hig
+ 2.174000000e-07 V_hig
+ 2.174010000e-07 V_hig
+ 2.175000000e-07 V_hig
+ 2.175010000e-07 V_hig
+ 2.176000000e-07 V_hig
+ 2.176010000e-07 V_hig
+ 2.177000000e-07 V_hig
+ 2.177010000e-07 V_hig
+ 2.178000000e-07 V_hig
+ 2.178010000e-07 V_hig
+ 2.179000000e-07 V_hig
+ 2.179010000e-07 V_low
+ 2.180000000e-07 V_low
+ 2.180010000e-07 V_low
+ 2.181000000e-07 V_low
+ 2.181010000e-07 V_low
+ 2.182000000e-07 V_low
+ 2.182010000e-07 V_low
+ 2.183000000e-07 V_low
+ 2.183010000e-07 V_low
+ 2.184000000e-07 V_low
+ 2.184010000e-07 V_low
+ 2.185000000e-07 V_low
+ 2.185010000e-07 V_low
+ 2.186000000e-07 V_low
+ 2.186010000e-07 V_low
+ 2.187000000e-07 V_low
+ 2.187010000e-07 V_low
+ 2.188000000e-07 V_low
+ 2.188010000e-07 V_low
+ 2.189000000e-07 V_low
+ 2.189010000e-07 V_hig
+ 2.190000000e-07 V_hig
+ 2.190010000e-07 V_hig
+ 2.191000000e-07 V_hig
+ 2.191010000e-07 V_hig
+ 2.192000000e-07 V_hig
+ 2.192010000e-07 V_hig
+ 2.193000000e-07 V_hig
+ 2.193010000e-07 V_hig
+ 2.194000000e-07 V_hig
+ 2.194010000e-07 V_hig
+ 2.195000000e-07 V_hig
+ 2.195010000e-07 V_hig
+ 2.196000000e-07 V_hig
+ 2.196010000e-07 V_hig
+ 2.197000000e-07 V_hig
+ 2.197010000e-07 V_hig
+ 2.198000000e-07 V_hig
+ 2.198010000e-07 V_hig
+ 2.199000000e-07 V_hig
+ 2.199010000e-07 V_hig
+ 2.200000000e-07 V_hig
+ 2.200010000e-07 V_hig
+ 2.201000000e-07 V_hig
+ 2.201010000e-07 V_hig
+ 2.202000000e-07 V_hig
+ 2.202010000e-07 V_hig
+ 2.203000000e-07 V_hig
+ 2.203010000e-07 V_hig
+ 2.204000000e-07 V_hig
+ 2.204010000e-07 V_hig
+ 2.205000000e-07 V_hig
+ 2.205010000e-07 V_hig
+ 2.206000000e-07 V_hig
+ 2.206010000e-07 V_hig
+ 2.207000000e-07 V_hig
+ 2.207010000e-07 V_hig
+ 2.208000000e-07 V_hig
+ 2.208010000e-07 V_hig
+ 2.209000000e-07 V_hig
+ 2.209010000e-07 V_low
+ 2.210000000e-07 V_low
+ 2.210010000e-07 V_low
+ 2.211000000e-07 V_low
+ 2.211010000e-07 V_low
+ 2.212000000e-07 V_low
+ 2.212010000e-07 V_low
+ 2.213000000e-07 V_low
+ 2.213010000e-07 V_low
+ 2.214000000e-07 V_low
+ 2.214010000e-07 V_low
+ 2.215000000e-07 V_low
+ 2.215010000e-07 V_low
+ 2.216000000e-07 V_low
+ 2.216010000e-07 V_low
+ 2.217000000e-07 V_low
+ 2.217010000e-07 V_low
+ 2.218000000e-07 V_low
+ 2.218010000e-07 V_low
+ 2.219000000e-07 V_low
+ 2.219010000e-07 V_low
+ 2.220000000e-07 V_low
+ 2.220010000e-07 V_low
+ 2.221000000e-07 V_low
+ 2.221010000e-07 V_low
+ 2.222000000e-07 V_low
+ 2.222010000e-07 V_low
+ 2.223000000e-07 V_low
+ 2.223010000e-07 V_low
+ 2.224000000e-07 V_low
+ 2.224010000e-07 V_low
+ 2.225000000e-07 V_low
+ 2.225010000e-07 V_low
+ 2.226000000e-07 V_low
+ 2.226010000e-07 V_low
+ 2.227000000e-07 V_low
+ 2.227010000e-07 V_low
+ 2.228000000e-07 V_low
+ 2.228010000e-07 V_low
+ 2.229000000e-07 V_low
+ 2.229010000e-07 V_hig
+ 2.230000000e-07 V_hig
+ 2.230010000e-07 V_hig
+ 2.231000000e-07 V_hig
+ 2.231010000e-07 V_hig
+ 2.232000000e-07 V_hig
+ 2.232010000e-07 V_hig
+ 2.233000000e-07 V_hig
+ 2.233010000e-07 V_hig
+ 2.234000000e-07 V_hig
+ 2.234010000e-07 V_hig
+ 2.235000000e-07 V_hig
+ 2.235010000e-07 V_hig
+ 2.236000000e-07 V_hig
+ 2.236010000e-07 V_hig
+ 2.237000000e-07 V_hig
+ 2.237010000e-07 V_hig
+ 2.238000000e-07 V_hig
+ 2.238010000e-07 V_hig
+ 2.239000000e-07 V_hig
+ 2.239010000e-07 V_hig
+ 2.240000000e-07 V_hig
+ 2.240010000e-07 V_hig
+ 2.241000000e-07 V_hig
+ 2.241010000e-07 V_hig
+ 2.242000000e-07 V_hig
+ 2.242010000e-07 V_hig
+ 2.243000000e-07 V_hig
+ 2.243010000e-07 V_hig
+ 2.244000000e-07 V_hig
+ 2.244010000e-07 V_hig
+ 2.245000000e-07 V_hig
+ 2.245010000e-07 V_hig
+ 2.246000000e-07 V_hig
+ 2.246010000e-07 V_hig
+ 2.247000000e-07 V_hig
+ 2.247010000e-07 V_hig
+ 2.248000000e-07 V_hig
+ 2.248010000e-07 V_hig
+ 2.249000000e-07 V_hig
+ 2.249010000e-07 V_hig
+ 2.250000000e-07 V_hig
+ 2.250010000e-07 V_hig
+ 2.251000000e-07 V_hig
+ 2.251010000e-07 V_hig
+ 2.252000000e-07 V_hig
+ 2.252010000e-07 V_hig
+ 2.253000000e-07 V_hig
+ 2.253010000e-07 V_hig
+ 2.254000000e-07 V_hig
+ 2.254010000e-07 V_hig
+ 2.255000000e-07 V_hig
+ 2.255010000e-07 V_hig
+ 2.256000000e-07 V_hig
+ 2.256010000e-07 V_hig
+ 2.257000000e-07 V_hig
+ 2.257010000e-07 V_hig
+ 2.258000000e-07 V_hig
+ 2.258010000e-07 V_hig
+ 2.259000000e-07 V_hig
+ 2.259010000e-07 V_hig
+ 2.260000000e-07 V_hig
+ 2.260010000e-07 V_hig
+ 2.261000000e-07 V_hig
+ 2.261010000e-07 V_hig
+ 2.262000000e-07 V_hig
+ 2.262010000e-07 V_hig
+ 2.263000000e-07 V_hig
+ 2.263010000e-07 V_hig
+ 2.264000000e-07 V_hig
+ 2.264010000e-07 V_hig
+ 2.265000000e-07 V_hig
+ 2.265010000e-07 V_hig
+ 2.266000000e-07 V_hig
+ 2.266010000e-07 V_hig
+ 2.267000000e-07 V_hig
+ 2.267010000e-07 V_hig
+ 2.268000000e-07 V_hig
+ 2.268010000e-07 V_hig
+ 2.269000000e-07 V_hig
+ 2.269010000e-07 V_hig
+ 2.270000000e-07 V_hig
+ 2.270010000e-07 V_hig
+ 2.271000000e-07 V_hig
+ 2.271010000e-07 V_hig
+ 2.272000000e-07 V_hig
+ 2.272010000e-07 V_hig
+ 2.273000000e-07 V_hig
+ 2.273010000e-07 V_hig
+ 2.274000000e-07 V_hig
+ 2.274010000e-07 V_hig
+ 2.275000000e-07 V_hig
+ 2.275010000e-07 V_hig
+ 2.276000000e-07 V_hig
+ 2.276010000e-07 V_hig
+ 2.277000000e-07 V_hig
+ 2.277010000e-07 V_hig
+ 2.278000000e-07 V_hig
+ 2.278010000e-07 V_hig
+ 2.279000000e-07 V_hig
+ 2.279010000e-07 V_low
+ 2.280000000e-07 V_low
+ 2.280010000e-07 V_low
+ 2.281000000e-07 V_low
+ 2.281010000e-07 V_low
+ 2.282000000e-07 V_low
+ 2.282010000e-07 V_low
+ 2.283000000e-07 V_low
+ 2.283010000e-07 V_low
+ 2.284000000e-07 V_low
+ 2.284010000e-07 V_low
+ 2.285000000e-07 V_low
+ 2.285010000e-07 V_low
+ 2.286000000e-07 V_low
+ 2.286010000e-07 V_low
+ 2.287000000e-07 V_low
+ 2.287010000e-07 V_low
+ 2.288000000e-07 V_low
+ 2.288010000e-07 V_low
+ 2.289000000e-07 V_low
+ 2.289010000e-07 V_low
+ 2.290000000e-07 V_low
+ 2.290010000e-07 V_low
+ 2.291000000e-07 V_low
+ 2.291010000e-07 V_low
+ 2.292000000e-07 V_low
+ 2.292010000e-07 V_low
+ 2.293000000e-07 V_low
+ 2.293010000e-07 V_low
+ 2.294000000e-07 V_low
+ 2.294010000e-07 V_low
+ 2.295000000e-07 V_low
+ 2.295010000e-07 V_low
+ 2.296000000e-07 V_low
+ 2.296010000e-07 V_low
+ 2.297000000e-07 V_low
+ 2.297010000e-07 V_low
+ 2.298000000e-07 V_low
+ 2.298010000e-07 V_low
+ 2.299000000e-07 V_low
+ 2.299010000e-07 V_low
+ 2.300000000e-07 V_low
+ 2.300010000e-07 V_low
+ 2.301000000e-07 V_low
+ 2.301010000e-07 V_low
+ 2.302000000e-07 V_low
+ 2.302010000e-07 V_low
+ 2.303000000e-07 V_low
+ 2.303010000e-07 V_low
+ 2.304000000e-07 V_low
+ 2.304010000e-07 V_low
+ 2.305000000e-07 V_low
+ 2.305010000e-07 V_low
+ 2.306000000e-07 V_low
+ 2.306010000e-07 V_low
+ 2.307000000e-07 V_low
+ 2.307010000e-07 V_low
+ 2.308000000e-07 V_low
+ 2.308010000e-07 V_low
+ 2.309000000e-07 V_low
+ 2.309010000e-07 V_low
+ 2.310000000e-07 V_low
+ 2.310010000e-07 V_low
+ 2.311000000e-07 V_low
+ 2.311010000e-07 V_low
+ 2.312000000e-07 V_low
+ 2.312010000e-07 V_low
+ 2.313000000e-07 V_low
+ 2.313010000e-07 V_low
+ 2.314000000e-07 V_low
+ 2.314010000e-07 V_low
+ 2.315000000e-07 V_low
+ 2.315010000e-07 V_low
+ 2.316000000e-07 V_low
+ 2.316010000e-07 V_low
+ 2.317000000e-07 V_low
+ 2.317010000e-07 V_low
+ 2.318000000e-07 V_low
+ 2.318010000e-07 V_low
+ 2.319000000e-07 V_low
+ 2.319010000e-07 V_low
+ 2.320000000e-07 V_low
+ 2.320010000e-07 V_low
+ 2.321000000e-07 V_low
+ 2.321010000e-07 V_low
+ 2.322000000e-07 V_low
+ 2.322010000e-07 V_low
+ 2.323000000e-07 V_low
+ 2.323010000e-07 V_low
+ 2.324000000e-07 V_low
+ 2.324010000e-07 V_low
+ 2.325000000e-07 V_low
+ 2.325010000e-07 V_low
+ 2.326000000e-07 V_low
+ 2.326010000e-07 V_low
+ 2.327000000e-07 V_low
+ 2.327010000e-07 V_low
+ 2.328000000e-07 V_low
+ 2.328010000e-07 V_low
+ 2.329000000e-07 V_low
+ 2.329010000e-07 V_low
+ 2.330000000e-07 V_low
+ 2.330010000e-07 V_low
+ 2.331000000e-07 V_low
+ 2.331010000e-07 V_low
+ 2.332000000e-07 V_low
+ 2.332010000e-07 V_low
+ 2.333000000e-07 V_low
+ 2.333010000e-07 V_low
+ 2.334000000e-07 V_low
+ 2.334010000e-07 V_low
+ 2.335000000e-07 V_low
+ 2.335010000e-07 V_low
+ 2.336000000e-07 V_low
+ 2.336010000e-07 V_low
+ 2.337000000e-07 V_low
+ 2.337010000e-07 V_low
+ 2.338000000e-07 V_low
+ 2.338010000e-07 V_low
+ 2.339000000e-07 V_low
+ 2.339010000e-07 V_low
+ 2.340000000e-07 V_low
+ 2.340010000e-07 V_low
+ 2.341000000e-07 V_low
+ 2.341010000e-07 V_low
+ 2.342000000e-07 V_low
+ 2.342010000e-07 V_low
+ 2.343000000e-07 V_low
+ 2.343010000e-07 V_low
+ 2.344000000e-07 V_low
+ 2.344010000e-07 V_low
+ 2.345000000e-07 V_low
+ 2.345010000e-07 V_low
+ 2.346000000e-07 V_low
+ 2.346010000e-07 V_low
+ 2.347000000e-07 V_low
+ 2.347010000e-07 V_low
+ 2.348000000e-07 V_low
+ 2.348010000e-07 V_low
+ 2.349000000e-07 V_low
+ 2.349010000e-07 V_hig
+ 2.350000000e-07 V_hig
+ 2.350010000e-07 V_hig
+ 2.351000000e-07 V_hig
+ 2.351010000e-07 V_hig
+ 2.352000000e-07 V_hig
+ 2.352010000e-07 V_hig
+ 2.353000000e-07 V_hig
+ 2.353010000e-07 V_hig
+ 2.354000000e-07 V_hig
+ 2.354010000e-07 V_hig
+ 2.355000000e-07 V_hig
+ 2.355010000e-07 V_hig
+ 2.356000000e-07 V_hig
+ 2.356010000e-07 V_hig
+ 2.357000000e-07 V_hig
+ 2.357010000e-07 V_hig
+ 2.358000000e-07 V_hig
+ 2.358010000e-07 V_hig
+ 2.359000000e-07 V_hig
+ 2.359010000e-07 V_low
+ 2.360000000e-07 V_low
+ 2.360010000e-07 V_low
+ 2.361000000e-07 V_low
+ 2.361010000e-07 V_low
+ 2.362000000e-07 V_low
+ 2.362010000e-07 V_low
+ 2.363000000e-07 V_low
+ 2.363010000e-07 V_low
+ 2.364000000e-07 V_low
+ 2.364010000e-07 V_low
+ 2.365000000e-07 V_low
+ 2.365010000e-07 V_low
+ 2.366000000e-07 V_low
+ 2.366010000e-07 V_low
+ 2.367000000e-07 V_low
+ 2.367010000e-07 V_low
+ 2.368000000e-07 V_low
+ 2.368010000e-07 V_low
+ 2.369000000e-07 V_low
+ 2.369010000e-07 V_hig
+ 2.370000000e-07 V_hig
+ 2.370010000e-07 V_hig
+ 2.371000000e-07 V_hig
+ 2.371010000e-07 V_hig
+ 2.372000000e-07 V_hig
+ 2.372010000e-07 V_hig
+ 2.373000000e-07 V_hig
+ 2.373010000e-07 V_hig
+ 2.374000000e-07 V_hig
+ 2.374010000e-07 V_hig
+ 2.375000000e-07 V_hig
+ 2.375010000e-07 V_hig
+ 2.376000000e-07 V_hig
+ 2.376010000e-07 V_hig
+ 2.377000000e-07 V_hig
+ 2.377010000e-07 V_hig
+ 2.378000000e-07 V_hig
+ 2.378010000e-07 V_hig
+ 2.379000000e-07 V_hig
+ 2.379010000e-07 V_low
+ 2.380000000e-07 V_low
+ 2.380010000e-07 V_low
+ 2.381000000e-07 V_low
+ 2.381010000e-07 V_low
+ 2.382000000e-07 V_low
+ 2.382010000e-07 V_low
+ 2.383000000e-07 V_low
+ 2.383010000e-07 V_low
+ 2.384000000e-07 V_low
+ 2.384010000e-07 V_low
+ 2.385000000e-07 V_low
+ 2.385010000e-07 V_low
+ 2.386000000e-07 V_low
+ 2.386010000e-07 V_low
+ 2.387000000e-07 V_low
+ 2.387010000e-07 V_low
+ 2.388000000e-07 V_low
+ 2.388010000e-07 V_low
+ 2.389000000e-07 V_low
+ 2.389010000e-07 V_hig
+ 2.390000000e-07 V_hig
+ 2.390010000e-07 V_hig
+ 2.391000000e-07 V_hig
+ 2.391010000e-07 V_hig
+ 2.392000000e-07 V_hig
+ 2.392010000e-07 V_hig
+ 2.393000000e-07 V_hig
+ 2.393010000e-07 V_hig
+ 2.394000000e-07 V_hig
+ 2.394010000e-07 V_hig
+ 2.395000000e-07 V_hig
+ 2.395010000e-07 V_hig
+ 2.396000000e-07 V_hig
+ 2.396010000e-07 V_hig
+ 2.397000000e-07 V_hig
+ 2.397010000e-07 V_hig
+ 2.398000000e-07 V_hig
+ 2.398010000e-07 V_hig
+ 2.399000000e-07 V_hig
+ 2.399010000e-07 V_low
+ 2.400000000e-07 V_low
+ 2.400010000e-07 V_low
+ 2.401000000e-07 V_low
+ 2.401010000e-07 V_low
+ 2.402000000e-07 V_low
+ 2.402010000e-07 V_low
+ 2.403000000e-07 V_low
+ 2.403010000e-07 V_low
+ 2.404000000e-07 V_low
+ 2.404010000e-07 V_low
+ 2.405000000e-07 V_low
+ 2.405010000e-07 V_low
+ 2.406000000e-07 V_low
+ 2.406010000e-07 V_low
+ 2.407000000e-07 V_low
+ 2.407010000e-07 V_low
+ 2.408000000e-07 V_low
+ 2.408010000e-07 V_low
+ 2.409000000e-07 V_low
+ 2.409010000e-07 V_hig
+ 2.410000000e-07 V_hig
+ 2.410010000e-07 V_hig
+ 2.411000000e-07 V_hig
+ 2.411010000e-07 V_hig
+ 2.412000000e-07 V_hig
+ 2.412010000e-07 V_hig
+ 2.413000000e-07 V_hig
+ 2.413010000e-07 V_hig
+ 2.414000000e-07 V_hig
+ 2.414010000e-07 V_hig
+ 2.415000000e-07 V_hig
+ 2.415010000e-07 V_hig
+ 2.416000000e-07 V_hig
+ 2.416010000e-07 V_hig
+ 2.417000000e-07 V_hig
+ 2.417010000e-07 V_hig
+ 2.418000000e-07 V_hig
+ 2.418010000e-07 V_hig
+ 2.419000000e-07 V_hig
+ 2.419010000e-07 V_hig
+ 2.420000000e-07 V_hig
+ 2.420010000e-07 V_hig
+ 2.421000000e-07 V_hig
+ 2.421010000e-07 V_hig
+ 2.422000000e-07 V_hig
+ 2.422010000e-07 V_hig
+ 2.423000000e-07 V_hig
+ 2.423010000e-07 V_hig
+ 2.424000000e-07 V_hig
+ 2.424010000e-07 V_hig
+ 2.425000000e-07 V_hig
+ 2.425010000e-07 V_hig
+ 2.426000000e-07 V_hig
+ 2.426010000e-07 V_hig
+ 2.427000000e-07 V_hig
+ 2.427010000e-07 V_hig
+ 2.428000000e-07 V_hig
+ 2.428010000e-07 V_hig
+ 2.429000000e-07 V_hig
+ 2.429010000e-07 V_hig
+ 2.430000000e-07 V_hig
+ 2.430010000e-07 V_hig
+ 2.431000000e-07 V_hig
+ 2.431010000e-07 V_hig
+ 2.432000000e-07 V_hig
+ 2.432010000e-07 V_hig
+ 2.433000000e-07 V_hig
+ 2.433010000e-07 V_hig
+ 2.434000000e-07 V_hig
+ 2.434010000e-07 V_hig
+ 2.435000000e-07 V_hig
+ 2.435010000e-07 V_hig
+ 2.436000000e-07 V_hig
+ 2.436010000e-07 V_hig
+ 2.437000000e-07 V_hig
+ 2.437010000e-07 V_hig
+ 2.438000000e-07 V_hig
+ 2.438010000e-07 V_hig
+ 2.439000000e-07 V_hig
+ 2.439010000e-07 V_hig
+ 2.440000000e-07 V_hig
+ 2.440010000e-07 V_hig
+ 2.441000000e-07 V_hig
+ 2.441010000e-07 V_hig
+ 2.442000000e-07 V_hig
+ 2.442010000e-07 V_hig
+ 2.443000000e-07 V_hig
+ 2.443010000e-07 V_hig
+ 2.444000000e-07 V_hig
+ 2.444010000e-07 V_hig
+ 2.445000000e-07 V_hig
+ 2.445010000e-07 V_hig
+ 2.446000000e-07 V_hig
+ 2.446010000e-07 V_hig
+ 2.447000000e-07 V_hig
+ 2.447010000e-07 V_hig
+ 2.448000000e-07 V_hig
+ 2.448010000e-07 V_hig
+ 2.449000000e-07 V_hig
+ 2.449010000e-07 V_low
+ 2.450000000e-07 V_low
+ 2.450010000e-07 V_low
+ 2.451000000e-07 V_low
+ 2.451010000e-07 V_low
+ 2.452000000e-07 V_low
+ 2.452010000e-07 V_low
+ 2.453000000e-07 V_low
+ 2.453010000e-07 V_low
+ 2.454000000e-07 V_low
+ 2.454010000e-07 V_low
+ 2.455000000e-07 V_low
+ 2.455010000e-07 V_low
+ 2.456000000e-07 V_low
+ 2.456010000e-07 V_low
+ 2.457000000e-07 V_low
+ 2.457010000e-07 V_low
+ 2.458000000e-07 V_low
+ 2.458010000e-07 V_low
+ 2.459000000e-07 V_low
+ 2.459010000e-07 V_hig
+ 2.460000000e-07 V_hig
+ 2.460010000e-07 V_hig
+ 2.461000000e-07 V_hig
+ 2.461010000e-07 V_hig
+ 2.462000000e-07 V_hig
+ 2.462010000e-07 V_hig
+ 2.463000000e-07 V_hig
+ 2.463010000e-07 V_hig
+ 2.464000000e-07 V_hig
+ 2.464010000e-07 V_hig
+ 2.465000000e-07 V_hig
+ 2.465010000e-07 V_hig
+ 2.466000000e-07 V_hig
+ 2.466010000e-07 V_hig
+ 2.467000000e-07 V_hig
+ 2.467010000e-07 V_hig
+ 2.468000000e-07 V_hig
+ 2.468010000e-07 V_hig
+ 2.469000000e-07 V_hig
+ 2.469010000e-07 V_hig
+ 2.470000000e-07 V_hig
+ 2.470010000e-07 V_hig
+ 2.471000000e-07 V_hig
+ 2.471010000e-07 V_hig
+ 2.472000000e-07 V_hig
+ 2.472010000e-07 V_hig
+ 2.473000000e-07 V_hig
+ 2.473010000e-07 V_hig
+ 2.474000000e-07 V_hig
+ 2.474010000e-07 V_hig
+ 2.475000000e-07 V_hig
+ 2.475010000e-07 V_hig
+ 2.476000000e-07 V_hig
+ 2.476010000e-07 V_hig
+ 2.477000000e-07 V_hig
+ 2.477010000e-07 V_hig
+ 2.478000000e-07 V_hig
+ 2.478010000e-07 V_hig
+ 2.479000000e-07 V_hig
+ 2.479010000e-07 V_low
+ 2.480000000e-07 V_low
+ 2.480010000e-07 V_low
+ 2.481000000e-07 V_low
+ 2.481010000e-07 V_low
+ 2.482000000e-07 V_low
+ 2.482010000e-07 V_low
+ 2.483000000e-07 V_low
+ 2.483010000e-07 V_low
+ 2.484000000e-07 V_low
+ 2.484010000e-07 V_low
+ 2.485000000e-07 V_low
+ 2.485010000e-07 V_low
+ 2.486000000e-07 V_low
+ 2.486010000e-07 V_low
+ 2.487000000e-07 V_low
+ 2.487010000e-07 V_low
+ 2.488000000e-07 V_low
+ 2.488010000e-07 V_low
+ 2.489000000e-07 V_low
+ 2.489010000e-07 V_low
+ 2.490000000e-07 V_low
+ 2.490010000e-07 V_low
+ 2.491000000e-07 V_low
+ 2.491010000e-07 V_low
+ 2.492000000e-07 V_low
+ 2.492010000e-07 V_low
+ 2.493000000e-07 V_low
+ 2.493010000e-07 V_low
+ 2.494000000e-07 V_low
+ 2.494010000e-07 V_low
+ 2.495000000e-07 V_low
+ 2.495010000e-07 V_low
+ 2.496000000e-07 V_low
+ 2.496010000e-07 V_low
+ 2.497000000e-07 V_low
+ 2.497010000e-07 V_low
+ 2.498000000e-07 V_low
+ 2.498010000e-07 V_low
+ 2.499000000e-07 V_low
+ 2.499010000e-07 V_low
+ 2.500000000e-07 V_low
+ 2.500010000e-07 V_low
+ 2.501000000e-07 V_low
+ 2.501010000e-07 V_low
+ 2.502000000e-07 V_low
+ 2.502010000e-07 V_low
+ 2.503000000e-07 V_low
+ 2.503010000e-07 V_low
+ 2.504000000e-07 V_low
+ 2.504010000e-07 V_low
+ 2.505000000e-07 V_low
+ 2.505010000e-07 V_low
+ 2.506000000e-07 V_low
+ 2.506010000e-07 V_low
+ 2.507000000e-07 V_low
+ 2.507010000e-07 V_low
+ 2.508000000e-07 V_low
+ 2.508010000e-07 V_low
+ 2.509000000e-07 V_low
+ 2.509010000e-07 V_hig
+ 2.510000000e-07 V_hig
+ 2.510010000e-07 V_hig
+ 2.511000000e-07 V_hig
+ 2.511010000e-07 V_hig
+ 2.512000000e-07 V_hig
+ 2.512010000e-07 V_hig
+ 2.513000000e-07 V_hig
+ 2.513010000e-07 V_hig
+ 2.514000000e-07 V_hig
+ 2.514010000e-07 V_hig
+ 2.515000000e-07 V_hig
+ 2.515010000e-07 V_hig
+ 2.516000000e-07 V_hig
+ 2.516010000e-07 V_hig
+ 2.517000000e-07 V_hig
+ 2.517010000e-07 V_hig
+ 2.518000000e-07 V_hig
+ 2.518010000e-07 V_hig
+ 2.519000000e-07 V_hig
+ 2.519010000e-07 V_hig
+ 2.520000000e-07 V_hig
+ 2.520010000e-07 V_hig
+ 2.521000000e-07 V_hig
+ 2.521010000e-07 V_hig
+ 2.522000000e-07 V_hig
+ 2.522010000e-07 V_hig
+ 2.523000000e-07 V_hig
+ 2.523010000e-07 V_hig
+ 2.524000000e-07 V_hig
+ 2.524010000e-07 V_hig
+ 2.525000000e-07 V_hig
+ 2.525010000e-07 V_hig
+ 2.526000000e-07 V_hig
+ 2.526010000e-07 V_hig
+ 2.527000000e-07 V_hig
+ 2.527010000e-07 V_hig
+ 2.528000000e-07 V_hig
+ 2.528010000e-07 V_hig
+ 2.529000000e-07 V_hig
+ 2.529010000e-07 V_low
+ 2.530000000e-07 V_low
+ 2.530010000e-07 V_low
+ 2.531000000e-07 V_low
+ 2.531010000e-07 V_low
+ 2.532000000e-07 V_low
+ 2.532010000e-07 V_low
+ 2.533000000e-07 V_low
+ 2.533010000e-07 V_low
+ 2.534000000e-07 V_low
+ 2.534010000e-07 V_low
+ 2.535000000e-07 V_low
+ 2.535010000e-07 V_low
+ 2.536000000e-07 V_low
+ 2.536010000e-07 V_low
+ 2.537000000e-07 V_low
+ 2.537010000e-07 V_low
+ 2.538000000e-07 V_low
+ 2.538010000e-07 V_low
+ 2.539000000e-07 V_low
+ 2.539010000e-07 V_hig
+ 2.540000000e-07 V_hig
+ 2.540010000e-07 V_hig
+ 2.541000000e-07 V_hig
+ 2.541010000e-07 V_hig
+ 2.542000000e-07 V_hig
+ 2.542010000e-07 V_hig
+ 2.543000000e-07 V_hig
+ 2.543010000e-07 V_hig
+ 2.544000000e-07 V_hig
+ 2.544010000e-07 V_hig
+ 2.545000000e-07 V_hig
+ 2.545010000e-07 V_hig
+ 2.546000000e-07 V_hig
+ 2.546010000e-07 V_hig
+ 2.547000000e-07 V_hig
+ 2.547010000e-07 V_hig
+ 2.548000000e-07 V_hig
+ 2.548010000e-07 V_hig
+ 2.549000000e-07 V_hig
+ 2.549010000e-07 V_low
+ 2.550000000e-07 V_low
+ 2.550010000e-07 V_low
+ 2.551000000e-07 V_low
+ 2.551010000e-07 V_low
+ 2.552000000e-07 V_low
+ 2.552010000e-07 V_low
+ 2.553000000e-07 V_low
+ 2.553010000e-07 V_low
+ 2.554000000e-07 V_low
+ 2.554010000e-07 V_low
+ 2.555000000e-07 V_low
+ 2.555010000e-07 V_low
+ 2.556000000e-07 V_low
+ 2.556010000e-07 V_low
+ 2.557000000e-07 V_low
+ 2.557010000e-07 V_low
+ 2.558000000e-07 V_low
+ 2.558010000e-07 V_low
+ 2.559000000e-07 V_low
+ 2.559010000e-07 V_low
+ 2.560000000e-07 V_low
+ 2.560010000e-07 V_low
+ 2.561000000e-07 V_low
+ 2.561010000e-07 V_low
+ 2.562000000e-07 V_low
+ 2.562010000e-07 V_low
+ 2.563000000e-07 V_low
+ 2.563010000e-07 V_low
+ 2.564000000e-07 V_low
+ 2.564010000e-07 V_low
+ 2.565000000e-07 V_low
+ 2.565010000e-07 V_low
+ 2.566000000e-07 V_low
+ 2.566010000e-07 V_low
+ 2.567000000e-07 V_low
+ 2.567010000e-07 V_low
+ 2.568000000e-07 V_low
+ 2.568010000e-07 V_low
+ 2.569000000e-07 V_low
+ 2.569010000e-07 V_low
+ 2.570000000e-07 V_low
+ 2.570010000e-07 V_low
+ 2.571000000e-07 V_low
+ 2.571010000e-07 V_low
+ 2.572000000e-07 V_low
+ 2.572010000e-07 V_low
+ 2.573000000e-07 V_low
+ 2.573010000e-07 V_low
+ 2.574000000e-07 V_low
+ 2.574010000e-07 V_low
+ 2.575000000e-07 V_low
+ 2.575010000e-07 V_low
+ 2.576000000e-07 V_low
+ 2.576010000e-07 V_low
+ 2.577000000e-07 V_low
+ 2.577010000e-07 V_low
+ 2.578000000e-07 V_low
+ 2.578010000e-07 V_low
+ 2.579000000e-07 V_low
+ 2.579010000e-07 V_low
+ 2.580000000e-07 V_low
+ 2.580010000e-07 V_low
+ 2.581000000e-07 V_low
+ 2.581010000e-07 V_low
+ 2.582000000e-07 V_low
+ 2.582010000e-07 V_low
+ 2.583000000e-07 V_low
+ 2.583010000e-07 V_low
+ 2.584000000e-07 V_low
+ 2.584010000e-07 V_low
+ 2.585000000e-07 V_low
+ 2.585010000e-07 V_low
+ 2.586000000e-07 V_low
+ 2.586010000e-07 V_low
+ 2.587000000e-07 V_low
+ 2.587010000e-07 V_low
+ 2.588000000e-07 V_low
+ 2.588010000e-07 V_low
+ 2.589000000e-07 V_low
+ 2.589010000e-07 V_low
+ 2.590000000e-07 V_low
+ 2.590010000e-07 V_low
+ 2.591000000e-07 V_low
+ 2.591010000e-07 V_low
+ 2.592000000e-07 V_low
+ 2.592010000e-07 V_low
+ 2.593000000e-07 V_low
+ 2.593010000e-07 V_low
+ 2.594000000e-07 V_low
+ 2.594010000e-07 V_low
+ 2.595000000e-07 V_low
+ 2.595010000e-07 V_low
+ 2.596000000e-07 V_low
+ 2.596010000e-07 V_low
+ 2.597000000e-07 V_low
+ 2.597010000e-07 V_low
+ 2.598000000e-07 V_low
+ 2.598010000e-07 V_low
+ 2.599000000e-07 V_low
+ 2.599010000e-07 V_hig
+ 2.600000000e-07 V_hig
+ 2.600010000e-07 V_hig
+ 2.601000000e-07 V_hig
+ 2.601010000e-07 V_hig
+ 2.602000000e-07 V_hig
+ 2.602010000e-07 V_hig
+ 2.603000000e-07 V_hig
+ 2.603010000e-07 V_hig
+ 2.604000000e-07 V_hig
+ 2.604010000e-07 V_hig
+ 2.605000000e-07 V_hig
+ 2.605010000e-07 V_hig
+ 2.606000000e-07 V_hig
+ 2.606010000e-07 V_hig
+ 2.607000000e-07 V_hig
+ 2.607010000e-07 V_hig
+ 2.608000000e-07 V_hig
+ 2.608010000e-07 V_hig
+ 2.609000000e-07 V_hig
+ 2.609010000e-07 V_low
+ 2.610000000e-07 V_low
+ 2.610010000e-07 V_low
+ 2.611000000e-07 V_low
+ 2.611010000e-07 V_low
+ 2.612000000e-07 V_low
+ 2.612010000e-07 V_low
+ 2.613000000e-07 V_low
+ 2.613010000e-07 V_low
+ 2.614000000e-07 V_low
+ 2.614010000e-07 V_low
+ 2.615000000e-07 V_low
+ 2.615010000e-07 V_low
+ 2.616000000e-07 V_low
+ 2.616010000e-07 V_low
+ 2.617000000e-07 V_low
+ 2.617010000e-07 V_low
+ 2.618000000e-07 V_low
+ 2.618010000e-07 V_low
+ 2.619000000e-07 V_low
+ 2.619010000e-07 V_low
+ 2.620000000e-07 V_low
+ 2.620010000e-07 V_low
+ 2.621000000e-07 V_low
+ 2.621010000e-07 V_low
+ 2.622000000e-07 V_low
+ 2.622010000e-07 V_low
+ 2.623000000e-07 V_low
+ 2.623010000e-07 V_low
+ 2.624000000e-07 V_low
+ 2.624010000e-07 V_low
+ 2.625000000e-07 V_low
+ 2.625010000e-07 V_low
+ 2.626000000e-07 V_low
+ 2.626010000e-07 V_low
+ 2.627000000e-07 V_low
+ 2.627010000e-07 V_low
+ 2.628000000e-07 V_low
+ 2.628010000e-07 V_low
+ 2.629000000e-07 V_low
+ 2.629010000e-07 V_low
+ 2.630000000e-07 V_low
+ 2.630010000e-07 V_low
+ 2.631000000e-07 V_low
+ 2.631010000e-07 V_low
+ 2.632000000e-07 V_low
+ 2.632010000e-07 V_low
+ 2.633000000e-07 V_low
+ 2.633010000e-07 V_low
+ 2.634000000e-07 V_low
+ 2.634010000e-07 V_low
+ 2.635000000e-07 V_low
+ 2.635010000e-07 V_low
+ 2.636000000e-07 V_low
+ 2.636010000e-07 V_low
+ 2.637000000e-07 V_low
+ 2.637010000e-07 V_low
+ 2.638000000e-07 V_low
+ 2.638010000e-07 V_low
+ 2.639000000e-07 V_low
+ 2.639010000e-07 V_low
+ 2.640000000e-07 V_low
+ 2.640010000e-07 V_low
+ 2.641000000e-07 V_low
+ 2.641010000e-07 V_low
+ 2.642000000e-07 V_low
+ 2.642010000e-07 V_low
+ 2.643000000e-07 V_low
+ 2.643010000e-07 V_low
+ 2.644000000e-07 V_low
+ 2.644010000e-07 V_low
+ 2.645000000e-07 V_low
+ 2.645010000e-07 V_low
+ 2.646000000e-07 V_low
+ 2.646010000e-07 V_low
+ 2.647000000e-07 V_low
+ 2.647010000e-07 V_low
+ 2.648000000e-07 V_low
+ 2.648010000e-07 V_low
+ 2.649000000e-07 V_low
+ 2.649010000e-07 V_low
+ 2.650000000e-07 V_low
+ 2.650010000e-07 V_low
+ 2.651000000e-07 V_low
+ 2.651010000e-07 V_low
+ 2.652000000e-07 V_low
+ 2.652010000e-07 V_low
+ 2.653000000e-07 V_low
+ 2.653010000e-07 V_low
+ 2.654000000e-07 V_low
+ 2.654010000e-07 V_low
+ 2.655000000e-07 V_low
+ 2.655010000e-07 V_low
+ 2.656000000e-07 V_low
+ 2.656010000e-07 V_low
+ 2.657000000e-07 V_low
+ 2.657010000e-07 V_low
+ 2.658000000e-07 V_low
+ 2.658010000e-07 V_low
+ 2.659000000e-07 V_low
+ 2.659010000e-07 V_low
+ 2.660000000e-07 V_low
+ 2.660010000e-07 V_low
+ 2.661000000e-07 V_low
+ 2.661010000e-07 V_low
+ 2.662000000e-07 V_low
+ 2.662010000e-07 V_low
+ 2.663000000e-07 V_low
+ 2.663010000e-07 V_low
+ 2.664000000e-07 V_low
+ 2.664010000e-07 V_low
+ 2.665000000e-07 V_low
+ 2.665010000e-07 V_low
+ 2.666000000e-07 V_low
+ 2.666010000e-07 V_low
+ 2.667000000e-07 V_low
+ 2.667010000e-07 V_low
+ 2.668000000e-07 V_low
+ 2.668010000e-07 V_low
+ 2.669000000e-07 V_low
+ 2.669010000e-07 V_hig
+ 2.670000000e-07 V_hig
+ 2.670010000e-07 V_hig
+ 2.671000000e-07 V_hig
+ 2.671010000e-07 V_hig
+ 2.672000000e-07 V_hig
+ 2.672010000e-07 V_hig
+ 2.673000000e-07 V_hig
+ 2.673010000e-07 V_hig
+ 2.674000000e-07 V_hig
+ 2.674010000e-07 V_hig
+ 2.675000000e-07 V_hig
+ 2.675010000e-07 V_hig
+ 2.676000000e-07 V_hig
+ 2.676010000e-07 V_hig
+ 2.677000000e-07 V_hig
+ 2.677010000e-07 V_hig
+ 2.678000000e-07 V_hig
+ 2.678010000e-07 V_hig
+ 2.679000000e-07 V_hig
+ 2.679010000e-07 V_hig
+ 2.680000000e-07 V_hig
+ 2.680010000e-07 V_hig
+ 2.681000000e-07 V_hig
+ 2.681010000e-07 V_hig
+ 2.682000000e-07 V_hig
+ 2.682010000e-07 V_hig
+ 2.683000000e-07 V_hig
+ 2.683010000e-07 V_hig
+ 2.684000000e-07 V_hig
+ 2.684010000e-07 V_hig
+ 2.685000000e-07 V_hig
+ 2.685010000e-07 V_hig
+ 2.686000000e-07 V_hig
+ 2.686010000e-07 V_hig
+ 2.687000000e-07 V_hig
+ 2.687010000e-07 V_hig
+ 2.688000000e-07 V_hig
+ 2.688010000e-07 V_hig
+ 2.689000000e-07 V_hig
+ 2.689010000e-07 V_hig
+ 2.690000000e-07 V_hig
+ 2.690010000e-07 V_hig
+ 2.691000000e-07 V_hig
+ 2.691010000e-07 V_hig
+ 2.692000000e-07 V_hig
+ 2.692010000e-07 V_hig
+ 2.693000000e-07 V_hig
+ 2.693010000e-07 V_hig
+ 2.694000000e-07 V_hig
+ 2.694010000e-07 V_hig
+ 2.695000000e-07 V_hig
+ 2.695010000e-07 V_hig
+ 2.696000000e-07 V_hig
+ 2.696010000e-07 V_hig
+ 2.697000000e-07 V_hig
+ 2.697010000e-07 V_hig
+ 2.698000000e-07 V_hig
+ 2.698010000e-07 V_hig
+ 2.699000000e-07 V_hig
+ 2.699010000e-07 V_hig
+ 2.700000000e-07 V_hig
+ 2.700010000e-07 V_hig
+ 2.701000000e-07 V_hig
+ 2.701010000e-07 V_hig
+ 2.702000000e-07 V_hig
+ 2.702010000e-07 V_hig
+ 2.703000000e-07 V_hig
+ 2.703010000e-07 V_hig
+ 2.704000000e-07 V_hig
+ 2.704010000e-07 V_hig
+ 2.705000000e-07 V_hig
+ 2.705010000e-07 V_hig
+ 2.706000000e-07 V_hig
+ 2.706010000e-07 V_hig
+ 2.707000000e-07 V_hig
+ 2.707010000e-07 V_hig
+ 2.708000000e-07 V_hig
+ 2.708010000e-07 V_hig
+ 2.709000000e-07 V_hig
+ 2.709010000e-07 V_low
+ 2.710000000e-07 V_low
+ 2.710010000e-07 V_low
+ 2.711000000e-07 V_low
+ 2.711010000e-07 V_low
+ 2.712000000e-07 V_low
+ 2.712010000e-07 V_low
+ 2.713000000e-07 V_low
+ 2.713010000e-07 V_low
+ 2.714000000e-07 V_low
+ 2.714010000e-07 V_low
+ 2.715000000e-07 V_low
+ 2.715010000e-07 V_low
+ 2.716000000e-07 V_low
+ 2.716010000e-07 V_low
+ 2.717000000e-07 V_low
+ 2.717010000e-07 V_low
+ 2.718000000e-07 V_low
+ 2.718010000e-07 V_low
+ 2.719000000e-07 V_low
+ 2.719010000e-07 V_hig
+ 2.720000000e-07 V_hig
+ 2.720010000e-07 V_hig
+ 2.721000000e-07 V_hig
+ 2.721010000e-07 V_hig
+ 2.722000000e-07 V_hig
+ 2.722010000e-07 V_hig
+ 2.723000000e-07 V_hig
+ 2.723010000e-07 V_hig
+ 2.724000000e-07 V_hig
+ 2.724010000e-07 V_hig
+ 2.725000000e-07 V_hig
+ 2.725010000e-07 V_hig
+ 2.726000000e-07 V_hig
+ 2.726010000e-07 V_hig
+ 2.727000000e-07 V_hig
+ 2.727010000e-07 V_hig
+ 2.728000000e-07 V_hig
+ 2.728010000e-07 V_hig
+ 2.729000000e-07 V_hig
+ 2.729010000e-07 V_hig
+ 2.730000000e-07 V_hig
+ 2.730010000e-07 V_hig
+ 2.731000000e-07 V_hig
+ 2.731010000e-07 V_hig
+ 2.732000000e-07 V_hig
+ 2.732010000e-07 V_hig
+ 2.733000000e-07 V_hig
+ 2.733010000e-07 V_hig
+ 2.734000000e-07 V_hig
+ 2.734010000e-07 V_hig
+ 2.735000000e-07 V_hig
+ 2.735010000e-07 V_hig
+ 2.736000000e-07 V_hig
+ 2.736010000e-07 V_hig
+ 2.737000000e-07 V_hig
+ 2.737010000e-07 V_hig
+ 2.738000000e-07 V_hig
+ 2.738010000e-07 V_hig
+ 2.739000000e-07 V_hig
+ 2.739010000e-07 V_hig
+ 2.740000000e-07 V_hig
+ 2.740010000e-07 V_hig
+ 2.741000000e-07 V_hig
+ 2.741010000e-07 V_hig
+ 2.742000000e-07 V_hig
+ 2.742010000e-07 V_hig
+ 2.743000000e-07 V_hig
+ 2.743010000e-07 V_hig
+ 2.744000000e-07 V_hig
+ 2.744010000e-07 V_hig
+ 2.745000000e-07 V_hig
+ 2.745010000e-07 V_hig
+ 2.746000000e-07 V_hig
+ 2.746010000e-07 V_hig
+ 2.747000000e-07 V_hig
+ 2.747010000e-07 V_hig
+ 2.748000000e-07 V_hig
+ 2.748010000e-07 V_hig
+ 2.749000000e-07 V_hig
+ 2.749010000e-07 V_hig
+ 2.750000000e-07 V_hig
+ 2.750010000e-07 V_hig
+ 2.751000000e-07 V_hig
+ 2.751010000e-07 V_hig
+ 2.752000000e-07 V_hig
+ 2.752010000e-07 V_hig
+ 2.753000000e-07 V_hig
+ 2.753010000e-07 V_hig
+ 2.754000000e-07 V_hig
+ 2.754010000e-07 V_hig
+ 2.755000000e-07 V_hig
+ 2.755010000e-07 V_hig
+ 2.756000000e-07 V_hig
+ 2.756010000e-07 V_hig
+ 2.757000000e-07 V_hig
+ 2.757010000e-07 V_hig
+ 2.758000000e-07 V_hig
+ 2.758010000e-07 V_hig
+ 2.759000000e-07 V_hig
+ 2.759010000e-07 V_low
+ 2.760000000e-07 V_low
+ 2.760010000e-07 V_low
+ 2.761000000e-07 V_low
+ 2.761010000e-07 V_low
+ 2.762000000e-07 V_low
+ 2.762010000e-07 V_low
+ 2.763000000e-07 V_low
+ 2.763010000e-07 V_low
+ 2.764000000e-07 V_low
+ 2.764010000e-07 V_low
+ 2.765000000e-07 V_low
+ 2.765010000e-07 V_low
+ 2.766000000e-07 V_low
+ 2.766010000e-07 V_low
+ 2.767000000e-07 V_low
+ 2.767010000e-07 V_low
+ 2.768000000e-07 V_low
+ 2.768010000e-07 V_low
+ 2.769000000e-07 V_low
+ 2.769010000e-07 V_hig
+ 2.770000000e-07 V_hig
+ 2.770010000e-07 V_hig
+ 2.771000000e-07 V_hig
+ 2.771010000e-07 V_hig
+ 2.772000000e-07 V_hig
+ 2.772010000e-07 V_hig
+ 2.773000000e-07 V_hig
+ 2.773010000e-07 V_hig
+ 2.774000000e-07 V_hig
+ 2.774010000e-07 V_hig
+ 2.775000000e-07 V_hig
+ 2.775010000e-07 V_hig
+ 2.776000000e-07 V_hig
+ 2.776010000e-07 V_hig
+ 2.777000000e-07 V_hig
+ 2.777010000e-07 V_hig
+ 2.778000000e-07 V_hig
+ 2.778010000e-07 V_hig
+ 2.779000000e-07 V_hig
+ 2.779010000e-07 V_low
+ 2.780000000e-07 V_low
+ 2.780010000e-07 V_low
+ 2.781000000e-07 V_low
+ 2.781010000e-07 V_low
+ 2.782000000e-07 V_low
+ 2.782010000e-07 V_low
+ 2.783000000e-07 V_low
+ 2.783010000e-07 V_low
+ 2.784000000e-07 V_low
+ 2.784010000e-07 V_low
+ 2.785000000e-07 V_low
+ 2.785010000e-07 V_low
+ 2.786000000e-07 V_low
+ 2.786010000e-07 V_low
+ 2.787000000e-07 V_low
+ 2.787010000e-07 V_low
+ 2.788000000e-07 V_low
+ 2.788010000e-07 V_low
+ 2.789000000e-07 V_low
+ 2.789010000e-07 V_hig
+ 2.790000000e-07 V_hig
+ 2.790010000e-07 V_hig
+ 2.791000000e-07 V_hig
+ 2.791010000e-07 V_hig
+ 2.792000000e-07 V_hig
+ 2.792010000e-07 V_hig
+ 2.793000000e-07 V_hig
+ 2.793010000e-07 V_hig
+ 2.794000000e-07 V_hig
+ 2.794010000e-07 V_hig
+ 2.795000000e-07 V_hig
+ 2.795010000e-07 V_hig
+ 2.796000000e-07 V_hig
+ 2.796010000e-07 V_hig
+ 2.797000000e-07 V_hig
+ 2.797010000e-07 V_hig
+ 2.798000000e-07 V_hig
+ 2.798010000e-07 V_hig
+ 2.799000000e-07 V_hig
+ 2.799010000e-07 V_low
+ 2.800000000e-07 V_low
+ 2.800010000e-07 V_low
+ 2.801000000e-07 V_low
+ 2.801010000e-07 V_low
+ 2.802000000e-07 V_low
+ 2.802010000e-07 V_low
+ 2.803000000e-07 V_low
+ 2.803010000e-07 V_low
+ 2.804000000e-07 V_low
+ 2.804010000e-07 V_low
+ 2.805000000e-07 V_low
+ 2.805010000e-07 V_low
+ 2.806000000e-07 V_low
+ 2.806010000e-07 V_low
+ 2.807000000e-07 V_low
+ 2.807010000e-07 V_low
+ 2.808000000e-07 V_low
+ 2.808010000e-07 V_low
+ 2.809000000e-07 V_low
+ 2.809010000e-07 V_low
+ 2.810000000e-07 V_low
+ 2.810010000e-07 V_low
+ 2.811000000e-07 V_low
+ 2.811010000e-07 V_low
+ 2.812000000e-07 V_low
+ 2.812010000e-07 V_low
+ 2.813000000e-07 V_low
+ 2.813010000e-07 V_low
+ 2.814000000e-07 V_low
+ 2.814010000e-07 V_low
+ 2.815000000e-07 V_low
+ 2.815010000e-07 V_low
+ 2.816000000e-07 V_low
+ 2.816010000e-07 V_low
+ 2.817000000e-07 V_low
+ 2.817010000e-07 V_low
+ 2.818000000e-07 V_low
+ 2.818010000e-07 V_low
+ 2.819000000e-07 V_low
+ 2.819010000e-07 V_low
+ 2.820000000e-07 V_low
+ 2.820010000e-07 V_low
+ 2.821000000e-07 V_low
+ 2.821010000e-07 V_low
+ 2.822000000e-07 V_low
+ 2.822010000e-07 V_low
+ 2.823000000e-07 V_low
+ 2.823010000e-07 V_low
+ 2.824000000e-07 V_low
+ 2.824010000e-07 V_low
+ 2.825000000e-07 V_low
+ 2.825010000e-07 V_low
+ 2.826000000e-07 V_low
+ 2.826010000e-07 V_low
+ 2.827000000e-07 V_low
+ 2.827010000e-07 V_low
+ 2.828000000e-07 V_low
+ 2.828010000e-07 V_low
+ 2.829000000e-07 V_low
+ 2.829010000e-07 V_hig
+ 2.830000000e-07 V_hig
+ 2.830010000e-07 V_hig
+ 2.831000000e-07 V_hig
+ 2.831010000e-07 V_hig
+ 2.832000000e-07 V_hig
+ 2.832010000e-07 V_hig
+ 2.833000000e-07 V_hig
+ 2.833010000e-07 V_hig
+ 2.834000000e-07 V_hig
+ 2.834010000e-07 V_hig
+ 2.835000000e-07 V_hig
+ 2.835010000e-07 V_hig
+ 2.836000000e-07 V_hig
+ 2.836010000e-07 V_hig
+ 2.837000000e-07 V_hig
+ 2.837010000e-07 V_hig
+ 2.838000000e-07 V_hig
+ 2.838010000e-07 V_hig
+ 2.839000000e-07 V_hig
+ 2.839010000e-07 V_low
+ 2.840000000e-07 V_low
+ 2.840010000e-07 V_low
+ 2.841000000e-07 V_low
+ 2.841010000e-07 V_low
+ 2.842000000e-07 V_low
+ 2.842010000e-07 V_low
+ 2.843000000e-07 V_low
+ 2.843010000e-07 V_low
+ 2.844000000e-07 V_low
+ 2.844010000e-07 V_low
+ 2.845000000e-07 V_low
+ 2.845010000e-07 V_low
+ 2.846000000e-07 V_low
+ 2.846010000e-07 V_low
+ 2.847000000e-07 V_low
+ 2.847010000e-07 V_low
+ 2.848000000e-07 V_low
+ 2.848010000e-07 V_low
+ 2.849000000e-07 V_low
+ 2.849010000e-07 V_hig
+ 2.850000000e-07 V_hig
+ 2.850010000e-07 V_hig
+ 2.851000000e-07 V_hig
+ 2.851010000e-07 V_hig
+ 2.852000000e-07 V_hig
+ 2.852010000e-07 V_hig
+ 2.853000000e-07 V_hig
+ 2.853010000e-07 V_hig
+ 2.854000000e-07 V_hig
+ 2.854010000e-07 V_hig
+ 2.855000000e-07 V_hig
+ 2.855010000e-07 V_hig
+ 2.856000000e-07 V_hig
+ 2.856010000e-07 V_hig
+ 2.857000000e-07 V_hig
+ 2.857010000e-07 V_hig
+ 2.858000000e-07 V_hig
+ 2.858010000e-07 V_hig
+ 2.859000000e-07 V_hig
+ 2.859010000e-07 V_low
+ 2.860000000e-07 V_low
+ 2.860010000e-07 V_low
+ 2.861000000e-07 V_low
+ 2.861010000e-07 V_low
+ 2.862000000e-07 V_low
+ 2.862010000e-07 V_low
+ 2.863000000e-07 V_low
+ 2.863010000e-07 V_low
+ 2.864000000e-07 V_low
+ 2.864010000e-07 V_low
+ 2.865000000e-07 V_low
+ 2.865010000e-07 V_low
+ 2.866000000e-07 V_low
+ 2.866010000e-07 V_low
+ 2.867000000e-07 V_low
+ 2.867010000e-07 V_low
+ 2.868000000e-07 V_low
+ 2.868010000e-07 V_low
+ 2.869000000e-07 V_low
+ 2.869010000e-07 V_low
+ 2.870000000e-07 V_low
+ 2.870010000e-07 V_low
+ 2.871000000e-07 V_low
+ 2.871010000e-07 V_low
+ 2.872000000e-07 V_low
+ 2.872010000e-07 V_low
+ 2.873000000e-07 V_low
+ 2.873010000e-07 V_low
+ 2.874000000e-07 V_low
+ 2.874010000e-07 V_low
+ 2.875000000e-07 V_low
+ 2.875010000e-07 V_low
+ 2.876000000e-07 V_low
+ 2.876010000e-07 V_low
+ 2.877000000e-07 V_low
+ 2.877010000e-07 V_low
+ 2.878000000e-07 V_low
+ 2.878010000e-07 V_low
+ 2.879000000e-07 V_low
+ 2.879010000e-07 V_hig
+ 2.880000000e-07 V_hig
+ 2.880010000e-07 V_hig
+ 2.881000000e-07 V_hig
+ 2.881010000e-07 V_hig
+ 2.882000000e-07 V_hig
+ 2.882010000e-07 V_hig
+ 2.883000000e-07 V_hig
+ 2.883010000e-07 V_hig
+ 2.884000000e-07 V_hig
+ 2.884010000e-07 V_hig
+ 2.885000000e-07 V_hig
+ 2.885010000e-07 V_hig
+ 2.886000000e-07 V_hig
+ 2.886010000e-07 V_hig
+ 2.887000000e-07 V_hig
+ 2.887010000e-07 V_hig
+ 2.888000000e-07 V_hig
+ 2.888010000e-07 V_hig
+ 2.889000000e-07 V_hig
+ 2.889010000e-07 V_low
+ 2.890000000e-07 V_low
+ 2.890010000e-07 V_low
+ 2.891000000e-07 V_low
+ 2.891010000e-07 V_low
+ 2.892000000e-07 V_low
+ 2.892010000e-07 V_low
+ 2.893000000e-07 V_low
+ 2.893010000e-07 V_low
+ 2.894000000e-07 V_low
+ 2.894010000e-07 V_low
+ 2.895000000e-07 V_low
+ 2.895010000e-07 V_low
+ 2.896000000e-07 V_low
+ 2.896010000e-07 V_low
+ 2.897000000e-07 V_low
+ 2.897010000e-07 V_low
+ 2.898000000e-07 V_low
+ 2.898010000e-07 V_low
+ 2.899000000e-07 V_low
+ 2.899010000e-07 V_low
+ 2.900000000e-07 V_low
+ 2.900010000e-07 V_low
+ 2.901000000e-07 V_low
+ 2.901010000e-07 V_low
+ 2.902000000e-07 V_low
+ 2.902010000e-07 V_low
+ 2.903000000e-07 V_low
+ 2.903010000e-07 V_low
+ 2.904000000e-07 V_low
+ 2.904010000e-07 V_low
+ 2.905000000e-07 V_low
+ 2.905010000e-07 V_low
+ 2.906000000e-07 V_low
+ 2.906010000e-07 V_low
+ 2.907000000e-07 V_low
+ 2.907010000e-07 V_low
+ 2.908000000e-07 V_low
+ 2.908010000e-07 V_low
+ 2.909000000e-07 V_low
+ 2.909010000e-07 V_low
+ 2.910000000e-07 V_low
+ 2.910010000e-07 V_low
+ 2.911000000e-07 V_low
+ 2.911010000e-07 V_low
+ 2.912000000e-07 V_low
+ 2.912010000e-07 V_low
+ 2.913000000e-07 V_low
+ 2.913010000e-07 V_low
+ 2.914000000e-07 V_low
+ 2.914010000e-07 V_low
+ 2.915000000e-07 V_low
+ 2.915010000e-07 V_low
+ 2.916000000e-07 V_low
+ 2.916010000e-07 V_low
+ 2.917000000e-07 V_low
+ 2.917010000e-07 V_low
+ 2.918000000e-07 V_low
+ 2.918010000e-07 V_low
+ 2.919000000e-07 V_low
+ 2.919010000e-07 V_hig
+ 2.920000000e-07 V_hig
+ 2.920010000e-07 V_hig
+ 2.921000000e-07 V_hig
+ 2.921010000e-07 V_hig
+ 2.922000000e-07 V_hig
+ 2.922010000e-07 V_hig
+ 2.923000000e-07 V_hig
+ 2.923010000e-07 V_hig
+ 2.924000000e-07 V_hig
+ 2.924010000e-07 V_hig
+ 2.925000000e-07 V_hig
+ 2.925010000e-07 V_hig
+ 2.926000000e-07 V_hig
+ 2.926010000e-07 V_hig
+ 2.927000000e-07 V_hig
+ 2.927010000e-07 V_hig
+ 2.928000000e-07 V_hig
+ 2.928010000e-07 V_hig
+ 2.929000000e-07 V_hig
+ 2.929010000e-07 V_low
+ 2.930000000e-07 V_low
+ 2.930010000e-07 V_low
+ 2.931000000e-07 V_low
+ 2.931010000e-07 V_low
+ 2.932000000e-07 V_low
+ 2.932010000e-07 V_low
+ 2.933000000e-07 V_low
+ 2.933010000e-07 V_low
+ 2.934000000e-07 V_low
+ 2.934010000e-07 V_low
+ 2.935000000e-07 V_low
+ 2.935010000e-07 V_low
+ 2.936000000e-07 V_low
+ 2.936010000e-07 V_low
+ 2.937000000e-07 V_low
+ 2.937010000e-07 V_low
+ 2.938000000e-07 V_low
+ 2.938010000e-07 V_low
+ 2.939000000e-07 V_low
+ 2.939010000e-07 V_low
+ 2.940000000e-07 V_low
+ 2.940010000e-07 V_low
+ 2.941000000e-07 V_low
+ 2.941010000e-07 V_low
+ 2.942000000e-07 V_low
+ 2.942010000e-07 V_low
+ 2.943000000e-07 V_low
+ 2.943010000e-07 V_low
+ 2.944000000e-07 V_low
+ 2.944010000e-07 V_low
+ 2.945000000e-07 V_low
+ 2.945010000e-07 V_low
+ 2.946000000e-07 V_low
+ 2.946010000e-07 V_low
+ 2.947000000e-07 V_low
+ 2.947010000e-07 V_low
+ 2.948000000e-07 V_low
+ 2.948010000e-07 V_low
+ 2.949000000e-07 V_low
+ 2.949010000e-07 V_hig
+ 2.950000000e-07 V_hig
+ 2.950010000e-07 V_hig
+ 2.951000000e-07 V_hig
+ 2.951010000e-07 V_hig
+ 2.952000000e-07 V_hig
+ 2.952010000e-07 V_hig
+ 2.953000000e-07 V_hig
+ 2.953010000e-07 V_hig
+ 2.954000000e-07 V_hig
+ 2.954010000e-07 V_hig
+ 2.955000000e-07 V_hig
+ 2.955010000e-07 V_hig
+ 2.956000000e-07 V_hig
+ 2.956010000e-07 V_hig
+ 2.957000000e-07 V_hig
+ 2.957010000e-07 V_hig
+ 2.958000000e-07 V_hig
+ 2.958010000e-07 V_hig
+ 2.959000000e-07 V_hig
+ 2.959010000e-07 V_hig
+ 2.960000000e-07 V_hig
+ 2.960010000e-07 V_hig
+ 2.961000000e-07 V_hig
+ 2.961010000e-07 V_hig
+ 2.962000000e-07 V_hig
+ 2.962010000e-07 V_hig
+ 2.963000000e-07 V_hig
+ 2.963010000e-07 V_hig
+ 2.964000000e-07 V_hig
+ 2.964010000e-07 V_hig
+ 2.965000000e-07 V_hig
+ 2.965010000e-07 V_hig
+ 2.966000000e-07 V_hig
+ 2.966010000e-07 V_hig
+ 2.967000000e-07 V_hig
+ 2.967010000e-07 V_hig
+ 2.968000000e-07 V_hig
+ 2.968010000e-07 V_hig
+ 2.969000000e-07 V_hig
+ 2.969010000e-07 V_low
+ 2.970000000e-07 V_low
+ 2.970010000e-07 V_low
+ 2.971000000e-07 V_low
+ 2.971010000e-07 V_low
+ 2.972000000e-07 V_low
+ 2.972010000e-07 V_low
+ 2.973000000e-07 V_low
+ 2.973010000e-07 V_low
+ 2.974000000e-07 V_low
+ 2.974010000e-07 V_low
+ 2.975000000e-07 V_low
+ 2.975010000e-07 V_low
+ 2.976000000e-07 V_low
+ 2.976010000e-07 V_low
+ 2.977000000e-07 V_low
+ 2.977010000e-07 V_low
+ 2.978000000e-07 V_low
+ 2.978010000e-07 V_low
+ 2.979000000e-07 V_low
+ 2.979010000e-07 V_hig
+ 2.980000000e-07 V_hig
+ 2.980010000e-07 V_hig
+ 2.981000000e-07 V_hig
+ 2.981010000e-07 V_hig
+ 2.982000000e-07 V_hig
+ 2.982010000e-07 V_hig
+ 2.983000000e-07 V_hig
+ 2.983010000e-07 V_hig
+ 2.984000000e-07 V_hig
+ 2.984010000e-07 V_hig
+ 2.985000000e-07 V_hig
+ 2.985010000e-07 V_hig
+ 2.986000000e-07 V_hig
+ 2.986010000e-07 V_hig
+ 2.987000000e-07 V_hig
+ 2.987010000e-07 V_hig
+ 2.988000000e-07 V_hig
+ 2.988010000e-07 V_hig
+ 2.989000000e-07 V_hig
+ 2.989010000e-07 V_hig
+ 2.990000000e-07 V_hig
+ 2.990010000e-07 V_hig
+ 2.991000000e-07 V_hig
+ 2.991010000e-07 V_hig
+ 2.992000000e-07 V_hig
+ 2.992010000e-07 V_hig
+ 2.993000000e-07 V_hig
+ 2.993010000e-07 V_hig
+ 2.994000000e-07 V_hig
+ 2.994010000e-07 V_hig
+ 2.995000000e-07 V_hig
+ 2.995010000e-07 V_hig
+ 2.996000000e-07 V_hig
+ 2.996010000e-07 V_hig
+ 2.997000000e-07 V_hig
+ 2.997010000e-07 V_hig
+ 2.998000000e-07 V_hig
+ 2.998010000e-07 V_hig
+ 2.999000000e-07 V_hig
+ 2.999010000e-07 V_low
+ 3.000000000e-07 V_low
+ 3.000010000e-07 V_low
+ 3.001000000e-07 V_low
+ 3.001010000e-07 V_low
+ 3.002000000e-07 V_low
+ 3.002010000e-07 V_low
+ 3.003000000e-07 V_low
+ 3.003010000e-07 V_low
+ 3.004000000e-07 V_low
+ 3.004010000e-07 V_low
+ 3.005000000e-07 V_low
+ 3.005010000e-07 V_low
+ 3.006000000e-07 V_low
+ 3.006010000e-07 V_low
+ 3.007000000e-07 V_low
+ 3.007010000e-07 V_low
+ 3.008000000e-07 V_low
+ 3.008010000e-07 V_low
+ 3.009000000e-07 V_low
+ 3.009010000e-07 V_hig
+ 3.010000000e-07 V_hig
+ 3.010010000e-07 V_hig
+ 3.011000000e-07 V_hig
+ 3.011010000e-07 V_hig
+ 3.012000000e-07 V_hig
+ 3.012010000e-07 V_hig
+ 3.013000000e-07 V_hig
+ 3.013010000e-07 V_hig
+ 3.014000000e-07 V_hig
+ 3.014010000e-07 V_hig
+ 3.015000000e-07 V_hig
+ 3.015010000e-07 V_hig
+ 3.016000000e-07 V_hig
+ 3.016010000e-07 V_hig
+ 3.017000000e-07 V_hig
+ 3.017010000e-07 V_hig
+ 3.018000000e-07 V_hig
+ 3.018010000e-07 V_hig
+ 3.019000000e-07 V_hig
+ 3.019010000e-07 V_hig
+ 3.020000000e-07 V_hig
+ 3.020010000e-07 V_hig
+ 3.021000000e-07 V_hig
+ 3.021010000e-07 V_hig
+ 3.022000000e-07 V_hig
+ 3.022010000e-07 V_hig
+ 3.023000000e-07 V_hig
+ 3.023010000e-07 V_hig
+ 3.024000000e-07 V_hig
+ 3.024010000e-07 V_hig
+ 3.025000000e-07 V_hig
+ 3.025010000e-07 V_hig
+ 3.026000000e-07 V_hig
+ 3.026010000e-07 V_hig
+ 3.027000000e-07 V_hig
+ 3.027010000e-07 V_hig
+ 3.028000000e-07 V_hig
+ 3.028010000e-07 V_hig
+ 3.029000000e-07 V_hig
+ 3.029010000e-07 V_hig
+ 3.030000000e-07 V_hig
+ 3.030010000e-07 V_hig
+ 3.031000000e-07 V_hig
+ 3.031010000e-07 V_hig
+ 3.032000000e-07 V_hig
+ 3.032010000e-07 V_hig
+ 3.033000000e-07 V_hig
+ 3.033010000e-07 V_hig
+ 3.034000000e-07 V_hig
+ 3.034010000e-07 V_hig
+ 3.035000000e-07 V_hig
+ 3.035010000e-07 V_hig
+ 3.036000000e-07 V_hig
+ 3.036010000e-07 V_hig
+ 3.037000000e-07 V_hig
+ 3.037010000e-07 V_hig
+ 3.038000000e-07 V_hig
+ 3.038010000e-07 V_hig
+ 3.039000000e-07 V_hig
+ 3.039010000e-07 V_hig
+ 3.040000000e-07 V_hig
+ 3.040010000e-07 V_hig
+ 3.041000000e-07 V_hig
+ 3.041010000e-07 V_hig
+ 3.042000000e-07 V_hig
+ 3.042010000e-07 V_hig
+ 3.043000000e-07 V_hig
+ 3.043010000e-07 V_hig
+ 3.044000000e-07 V_hig
+ 3.044010000e-07 V_hig
+ 3.045000000e-07 V_hig
+ 3.045010000e-07 V_hig
+ 3.046000000e-07 V_hig
+ 3.046010000e-07 V_hig
+ 3.047000000e-07 V_hig
+ 3.047010000e-07 V_hig
+ 3.048000000e-07 V_hig
+ 3.048010000e-07 V_hig
+ 3.049000000e-07 V_hig
+ 3.049010000e-07 V_hig
+ 3.050000000e-07 V_hig
+ 3.050010000e-07 V_hig
+ 3.051000000e-07 V_hig
+ 3.051010000e-07 V_hig
+ 3.052000000e-07 V_hig
+ 3.052010000e-07 V_hig
+ 3.053000000e-07 V_hig
+ 3.053010000e-07 V_hig
+ 3.054000000e-07 V_hig
+ 3.054010000e-07 V_hig
+ 3.055000000e-07 V_hig
+ 3.055010000e-07 V_hig
+ 3.056000000e-07 V_hig
+ 3.056010000e-07 V_hig
+ 3.057000000e-07 V_hig
+ 3.057010000e-07 V_hig
+ 3.058000000e-07 V_hig
+ 3.058010000e-07 V_hig
+ 3.059000000e-07 V_hig
+ 3.059010000e-07 V_hig
+ 3.060000000e-07 V_hig
+ 3.060010000e-07 V_hig
+ 3.061000000e-07 V_hig
+ 3.061010000e-07 V_hig
+ 3.062000000e-07 V_hig
+ 3.062010000e-07 V_hig
+ 3.063000000e-07 V_hig
+ 3.063010000e-07 V_hig
+ 3.064000000e-07 V_hig
+ 3.064010000e-07 V_hig
+ 3.065000000e-07 V_hig
+ 3.065010000e-07 V_hig
+ 3.066000000e-07 V_hig
+ 3.066010000e-07 V_hig
+ 3.067000000e-07 V_hig
+ 3.067010000e-07 V_hig
+ 3.068000000e-07 V_hig
+ 3.068010000e-07 V_hig
+ 3.069000000e-07 V_hig
+ 3.069010000e-07 V_hig
+ 3.070000000e-07 V_hig
+ 3.070010000e-07 V_hig
+ 3.071000000e-07 V_hig
+ 3.071010000e-07 V_hig
+ 3.072000000e-07 V_hig
+ 3.072010000e-07 V_hig
+ 3.073000000e-07 V_hig
+ 3.073010000e-07 V_hig
+ 3.074000000e-07 V_hig
+ 3.074010000e-07 V_hig
+ 3.075000000e-07 V_hig
+ 3.075010000e-07 V_hig
+ 3.076000000e-07 V_hig
+ 3.076010000e-07 V_hig
+ 3.077000000e-07 V_hig
+ 3.077010000e-07 V_hig
+ 3.078000000e-07 V_hig
+ 3.078010000e-07 V_hig
+ 3.079000000e-07 V_hig
+ 3.079010000e-07 V_low
+ 3.080000000e-07 V_low
+ 3.080010000e-07 V_low
+ 3.081000000e-07 V_low
+ 3.081010000e-07 V_low
+ 3.082000000e-07 V_low
+ 3.082010000e-07 V_low
+ 3.083000000e-07 V_low
+ 3.083010000e-07 V_low
+ 3.084000000e-07 V_low
+ 3.084010000e-07 V_low
+ 3.085000000e-07 V_low
+ 3.085010000e-07 V_low
+ 3.086000000e-07 V_low
+ 3.086010000e-07 V_low
+ 3.087000000e-07 V_low
+ 3.087010000e-07 V_low
+ 3.088000000e-07 V_low
+ 3.088010000e-07 V_low
+ 3.089000000e-07 V_low
+ 3.089010000e-07 V_low
+ 3.090000000e-07 V_low
+ 3.090010000e-07 V_low
+ 3.091000000e-07 V_low
+ 3.091010000e-07 V_low
+ 3.092000000e-07 V_low
+ 3.092010000e-07 V_low
+ 3.093000000e-07 V_low
+ 3.093010000e-07 V_low
+ 3.094000000e-07 V_low
+ 3.094010000e-07 V_low
+ 3.095000000e-07 V_low
+ 3.095010000e-07 V_low
+ 3.096000000e-07 V_low
+ 3.096010000e-07 V_low
+ 3.097000000e-07 V_low
+ 3.097010000e-07 V_low
+ 3.098000000e-07 V_low
+ 3.098010000e-07 V_low
+ 3.099000000e-07 V_low
+ 3.099010000e-07 V_low
+ 3.100000000e-07 V_low
+ 3.100010000e-07 V_low
+ 3.101000000e-07 V_low
+ 3.101010000e-07 V_low
+ 3.102000000e-07 V_low
+ 3.102010000e-07 V_low
+ 3.103000000e-07 V_low
+ 3.103010000e-07 V_low
+ 3.104000000e-07 V_low
+ 3.104010000e-07 V_low
+ 3.105000000e-07 V_low
+ 3.105010000e-07 V_low
+ 3.106000000e-07 V_low
+ 3.106010000e-07 V_low
+ 3.107000000e-07 V_low
+ 3.107010000e-07 V_low
+ 3.108000000e-07 V_low
+ 3.108010000e-07 V_low
+ 3.109000000e-07 V_low
+ 3.109010000e-07 V_low
+ 3.110000000e-07 V_low
+ 3.110010000e-07 V_low
+ 3.111000000e-07 V_low
+ 3.111010000e-07 V_low
+ 3.112000000e-07 V_low
+ 3.112010000e-07 V_low
+ 3.113000000e-07 V_low
+ 3.113010000e-07 V_low
+ 3.114000000e-07 V_low
+ 3.114010000e-07 V_low
+ 3.115000000e-07 V_low
+ 3.115010000e-07 V_low
+ 3.116000000e-07 V_low
+ 3.116010000e-07 V_low
+ 3.117000000e-07 V_low
+ 3.117010000e-07 V_low
+ 3.118000000e-07 V_low
+ 3.118010000e-07 V_low
+ 3.119000000e-07 V_low
+ 3.119010000e-07 V_hig
+ 3.120000000e-07 V_hig
+ 3.120010000e-07 V_hig
+ 3.121000000e-07 V_hig
+ 3.121010000e-07 V_hig
+ 3.122000000e-07 V_hig
+ 3.122010000e-07 V_hig
+ 3.123000000e-07 V_hig
+ 3.123010000e-07 V_hig
+ 3.124000000e-07 V_hig
+ 3.124010000e-07 V_hig
+ 3.125000000e-07 V_hig
+ 3.125010000e-07 V_hig
+ 3.126000000e-07 V_hig
+ 3.126010000e-07 V_hig
+ 3.127000000e-07 V_hig
+ 3.127010000e-07 V_hig
+ 3.128000000e-07 V_hig
+ 3.128010000e-07 V_hig
+ 3.129000000e-07 V_hig
+ 3.129010000e-07 V_hig
+ 3.130000000e-07 V_hig
+ 3.130010000e-07 V_hig
+ 3.131000000e-07 V_hig
+ 3.131010000e-07 V_hig
+ 3.132000000e-07 V_hig
+ 3.132010000e-07 V_hig
+ 3.133000000e-07 V_hig
+ 3.133010000e-07 V_hig
+ 3.134000000e-07 V_hig
+ 3.134010000e-07 V_hig
+ 3.135000000e-07 V_hig
+ 3.135010000e-07 V_hig
+ 3.136000000e-07 V_hig
+ 3.136010000e-07 V_hig
+ 3.137000000e-07 V_hig
+ 3.137010000e-07 V_hig
+ 3.138000000e-07 V_hig
+ 3.138010000e-07 V_hig
+ 3.139000000e-07 V_hig
+ 3.139010000e-07 V_low
+ 3.140000000e-07 V_low
+ 3.140010000e-07 V_low
+ 3.141000000e-07 V_low
+ 3.141010000e-07 V_low
+ 3.142000000e-07 V_low
+ 3.142010000e-07 V_low
+ 3.143000000e-07 V_low
+ 3.143010000e-07 V_low
+ 3.144000000e-07 V_low
+ 3.144010000e-07 V_low
+ 3.145000000e-07 V_low
+ 3.145010000e-07 V_low
+ 3.146000000e-07 V_low
+ 3.146010000e-07 V_low
+ 3.147000000e-07 V_low
+ 3.147010000e-07 V_low
+ 3.148000000e-07 V_low
+ 3.148010000e-07 V_low
+ 3.149000000e-07 V_low
+ 3.149010000e-07 V_low
+ 3.150000000e-07 V_low
+ 3.150010000e-07 V_low
+ 3.151000000e-07 V_low
+ 3.151010000e-07 V_low
+ 3.152000000e-07 V_low
+ 3.152010000e-07 V_low
+ 3.153000000e-07 V_low
+ 3.153010000e-07 V_low
+ 3.154000000e-07 V_low
+ 3.154010000e-07 V_low
+ 3.155000000e-07 V_low
+ 3.155010000e-07 V_low
+ 3.156000000e-07 V_low
+ 3.156010000e-07 V_low
+ 3.157000000e-07 V_low
+ 3.157010000e-07 V_low
+ 3.158000000e-07 V_low
+ 3.158010000e-07 V_low
+ 3.159000000e-07 V_low
+ 3.159010000e-07 V_hig
+ 3.160000000e-07 V_hig
+ 3.160010000e-07 V_hig
+ 3.161000000e-07 V_hig
+ 3.161010000e-07 V_hig
+ 3.162000000e-07 V_hig
+ 3.162010000e-07 V_hig
+ 3.163000000e-07 V_hig
+ 3.163010000e-07 V_hig
+ 3.164000000e-07 V_hig
+ 3.164010000e-07 V_hig
+ 3.165000000e-07 V_hig
+ 3.165010000e-07 V_hig
+ 3.166000000e-07 V_hig
+ 3.166010000e-07 V_hig
+ 3.167000000e-07 V_hig
+ 3.167010000e-07 V_hig
+ 3.168000000e-07 V_hig
+ 3.168010000e-07 V_hig
+ 3.169000000e-07 V_hig
+ 3.169010000e-07 V_hig
+ 3.170000000e-07 V_hig
+ 3.170010000e-07 V_hig
+ 3.171000000e-07 V_hig
+ 3.171010000e-07 V_hig
+ 3.172000000e-07 V_hig
+ 3.172010000e-07 V_hig
+ 3.173000000e-07 V_hig
+ 3.173010000e-07 V_hig
+ 3.174000000e-07 V_hig
+ 3.174010000e-07 V_hig
+ 3.175000000e-07 V_hig
+ 3.175010000e-07 V_hig
+ 3.176000000e-07 V_hig
+ 3.176010000e-07 V_hig
+ 3.177000000e-07 V_hig
+ 3.177010000e-07 V_hig
+ 3.178000000e-07 V_hig
+ 3.178010000e-07 V_hig
+ 3.179000000e-07 V_hig
+ 3.179010000e-07 V_hig
+ 3.180000000e-07 V_hig
+ 3.180010000e-07 V_hig
+ 3.181000000e-07 V_hig
+ 3.181010000e-07 V_hig
+ 3.182000000e-07 V_hig
+ 3.182010000e-07 V_hig
+ 3.183000000e-07 V_hig
+ 3.183010000e-07 V_hig
+ 3.184000000e-07 V_hig
+ 3.184010000e-07 V_hig
+ 3.185000000e-07 V_hig
+ 3.185010000e-07 V_hig
+ 3.186000000e-07 V_hig
+ 3.186010000e-07 V_hig
+ 3.187000000e-07 V_hig
+ 3.187010000e-07 V_hig
+ 3.188000000e-07 V_hig
+ 3.188010000e-07 V_hig
+ 3.189000000e-07 V_hig
+ 3.189010000e-07 V_hig
+ 3.190000000e-07 V_hig
+ 3.190010000e-07 V_hig
+ 3.191000000e-07 V_hig
+ 3.191010000e-07 V_hig
+ 3.192000000e-07 V_hig
+ 3.192010000e-07 V_hig
+ 3.193000000e-07 V_hig
+ 3.193010000e-07 V_hig
+ 3.194000000e-07 V_hig
+ 3.194010000e-07 V_hig
+ 3.195000000e-07 V_hig
+ 3.195010000e-07 V_hig
+ 3.196000000e-07 V_hig
+ 3.196010000e-07 V_hig
+ 3.197000000e-07 V_hig
+ 3.197010000e-07 V_hig
+ 3.198000000e-07 V_hig
+ 3.198010000e-07 V_hig
+ 3.199000000e-07 V_hig
+ 3.199010000e-07 V_hig
+ 3.200000000e-07 V_hig
+ 3.200010000e-07 V_hig
+ 3.201000000e-07 V_hig
+ 3.201010000e-07 V_hig
+ 3.202000000e-07 V_hig
+ 3.202010000e-07 V_hig
+ 3.203000000e-07 V_hig
+ 3.203010000e-07 V_hig
+ 3.204000000e-07 V_hig
+ 3.204010000e-07 V_hig
+ 3.205000000e-07 V_hig
+ 3.205010000e-07 V_hig
+ 3.206000000e-07 V_hig
+ 3.206010000e-07 V_hig
+ 3.207000000e-07 V_hig
+ 3.207010000e-07 V_hig
+ 3.208000000e-07 V_hig
+ 3.208010000e-07 V_hig
+ 3.209000000e-07 V_hig
+ 3.209010000e-07 V_hig
+ 3.210000000e-07 V_hig
+ 3.210010000e-07 V_hig
+ 3.211000000e-07 V_hig
+ 3.211010000e-07 V_hig
+ 3.212000000e-07 V_hig
+ 3.212010000e-07 V_hig
+ 3.213000000e-07 V_hig
+ 3.213010000e-07 V_hig
+ 3.214000000e-07 V_hig
+ 3.214010000e-07 V_hig
+ 3.215000000e-07 V_hig
+ 3.215010000e-07 V_hig
+ 3.216000000e-07 V_hig
+ 3.216010000e-07 V_hig
+ 3.217000000e-07 V_hig
+ 3.217010000e-07 V_hig
+ 3.218000000e-07 V_hig
+ 3.218010000e-07 V_hig
+ 3.219000000e-07 V_hig
+ 3.219010000e-07 V_hig
+ 3.220000000e-07 V_hig
+ 3.220010000e-07 V_hig
+ 3.221000000e-07 V_hig
+ 3.221010000e-07 V_hig
+ 3.222000000e-07 V_hig
+ 3.222010000e-07 V_hig
+ 3.223000000e-07 V_hig
+ 3.223010000e-07 V_hig
+ 3.224000000e-07 V_hig
+ 3.224010000e-07 V_hig
+ 3.225000000e-07 V_hig
+ 3.225010000e-07 V_hig
+ 3.226000000e-07 V_hig
+ 3.226010000e-07 V_hig
+ 3.227000000e-07 V_hig
+ 3.227010000e-07 V_hig
+ 3.228000000e-07 V_hig
+ 3.228010000e-07 V_hig
+ 3.229000000e-07 V_hig
+ 3.229010000e-07 V_low
+ 3.230000000e-07 V_low
+ 3.230010000e-07 V_low
+ 3.231000000e-07 V_low
+ 3.231010000e-07 V_low
+ 3.232000000e-07 V_low
+ 3.232010000e-07 V_low
+ 3.233000000e-07 V_low
+ 3.233010000e-07 V_low
+ 3.234000000e-07 V_low
+ 3.234010000e-07 V_low
+ 3.235000000e-07 V_low
+ 3.235010000e-07 V_low
+ 3.236000000e-07 V_low
+ 3.236010000e-07 V_low
+ 3.237000000e-07 V_low
+ 3.237010000e-07 V_low
+ 3.238000000e-07 V_low
+ 3.238010000e-07 V_low
+ 3.239000000e-07 V_low
+ 3.239010000e-07 V_hig
+ 3.240000000e-07 V_hig
+ 3.240010000e-07 V_hig
+ 3.241000000e-07 V_hig
+ 3.241010000e-07 V_hig
+ 3.242000000e-07 V_hig
+ 3.242010000e-07 V_hig
+ 3.243000000e-07 V_hig
+ 3.243010000e-07 V_hig
+ 3.244000000e-07 V_hig
+ 3.244010000e-07 V_hig
+ 3.245000000e-07 V_hig
+ 3.245010000e-07 V_hig
+ 3.246000000e-07 V_hig
+ 3.246010000e-07 V_hig
+ 3.247000000e-07 V_hig
+ 3.247010000e-07 V_hig
+ 3.248000000e-07 V_hig
+ 3.248010000e-07 V_hig
+ 3.249000000e-07 V_hig
+ 3.249010000e-07 V_low
+ 3.250000000e-07 V_low
+ 3.250010000e-07 V_low
+ 3.251000000e-07 V_low
+ 3.251010000e-07 V_low
+ 3.252000000e-07 V_low
+ 3.252010000e-07 V_low
+ 3.253000000e-07 V_low
+ 3.253010000e-07 V_low
+ 3.254000000e-07 V_low
+ 3.254010000e-07 V_low
+ 3.255000000e-07 V_low
+ 3.255010000e-07 V_low
+ 3.256000000e-07 V_low
+ 3.256010000e-07 V_low
+ 3.257000000e-07 V_low
+ 3.257010000e-07 V_low
+ 3.258000000e-07 V_low
+ 3.258010000e-07 V_low
+ 3.259000000e-07 V_low
+ 3.259010000e-07 V_low
+ 3.260000000e-07 V_low
+ 3.260010000e-07 V_low
+ 3.261000000e-07 V_low
+ 3.261010000e-07 V_low
+ 3.262000000e-07 V_low
+ 3.262010000e-07 V_low
+ 3.263000000e-07 V_low
+ 3.263010000e-07 V_low
+ 3.264000000e-07 V_low
+ 3.264010000e-07 V_low
+ 3.265000000e-07 V_low
+ 3.265010000e-07 V_low
+ 3.266000000e-07 V_low
+ 3.266010000e-07 V_low
+ 3.267000000e-07 V_low
+ 3.267010000e-07 V_low
+ 3.268000000e-07 V_low
+ 3.268010000e-07 V_low
+ 3.269000000e-07 V_low
+ 3.269010000e-07 V_hig
+ 3.270000000e-07 V_hig
+ 3.270010000e-07 V_hig
+ 3.271000000e-07 V_hig
+ 3.271010000e-07 V_hig
+ 3.272000000e-07 V_hig
+ 3.272010000e-07 V_hig
+ 3.273000000e-07 V_hig
+ 3.273010000e-07 V_hig
+ 3.274000000e-07 V_hig
+ 3.274010000e-07 V_hig
+ 3.275000000e-07 V_hig
+ 3.275010000e-07 V_hig
+ 3.276000000e-07 V_hig
+ 3.276010000e-07 V_hig
+ 3.277000000e-07 V_hig
+ 3.277010000e-07 V_hig
+ 3.278000000e-07 V_hig
+ 3.278010000e-07 V_hig
+ 3.279000000e-07 V_hig
+ 3.279010000e-07 V_hig
+ 3.280000000e-07 V_hig
+ 3.280010000e-07 V_hig
+ 3.281000000e-07 V_hig
+ 3.281010000e-07 V_hig
+ 3.282000000e-07 V_hig
+ 3.282010000e-07 V_hig
+ 3.283000000e-07 V_hig
+ 3.283010000e-07 V_hig
+ 3.284000000e-07 V_hig
+ 3.284010000e-07 V_hig
+ 3.285000000e-07 V_hig
+ 3.285010000e-07 V_hig
+ 3.286000000e-07 V_hig
+ 3.286010000e-07 V_hig
+ 3.287000000e-07 V_hig
+ 3.287010000e-07 V_hig
+ 3.288000000e-07 V_hig
+ 3.288010000e-07 V_hig
+ 3.289000000e-07 V_hig
+ 3.289010000e-07 V_low
+ 3.290000000e-07 V_low
+ 3.290010000e-07 V_low
+ 3.291000000e-07 V_low
+ 3.291010000e-07 V_low
+ 3.292000000e-07 V_low
+ 3.292010000e-07 V_low
+ 3.293000000e-07 V_low
+ 3.293010000e-07 V_low
+ 3.294000000e-07 V_low
+ 3.294010000e-07 V_low
+ 3.295000000e-07 V_low
+ 3.295010000e-07 V_low
+ 3.296000000e-07 V_low
+ 3.296010000e-07 V_low
+ 3.297000000e-07 V_low
+ 3.297010000e-07 V_low
+ 3.298000000e-07 V_low
+ 3.298010000e-07 V_low
+ 3.299000000e-07 V_low
+ 3.299010000e-07 V_hig
+ 3.300000000e-07 V_hig
+ 3.300010000e-07 V_hig
+ 3.301000000e-07 V_hig
+ 3.301010000e-07 V_hig
+ 3.302000000e-07 V_hig
+ 3.302010000e-07 V_hig
+ 3.303000000e-07 V_hig
+ 3.303010000e-07 V_hig
+ 3.304000000e-07 V_hig
+ 3.304010000e-07 V_hig
+ 3.305000000e-07 V_hig
+ 3.305010000e-07 V_hig
+ 3.306000000e-07 V_hig
+ 3.306010000e-07 V_hig
+ 3.307000000e-07 V_hig
+ 3.307010000e-07 V_hig
+ 3.308000000e-07 V_hig
+ 3.308010000e-07 V_hig
+ 3.309000000e-07 V_hig
+ 3.309010000e-07 V_hig
+ 3.310000000e-07 V_hig
+ 3.310010000e-07 V_hig
+ 3.311000000e-07 V_hig
+ 3.311010000e-07 V_hig
+ 3.312000000e-07 V_hig
+ 3.312010000e-07 V_hig
+ 3.313000000e-07 V_hig
+ 3.313010000e-07 V_hig
+ 3.314000000e-07 V_hig
+ 3.314010000e-07 V_hig
+ 3.315000000e-07 V_hig
+ 3.315010000e-07 V_hig
+ 3.316000000e-07 V_hig
+ 3.316010000e-07 V_hig
+ 3.317000000e-07 V_hig
+ 3.317010000e-07 V_hig
+ 3.318000000e-07 V_hig
+ 3.318010000e-07 V_hig
+ 3.319000000e-07 V_hig
+ 3.319010000e-07 V_hig
+ 3.320000000e-07 V_hig
+ 3.320010000e-07 V_hig
+ 3.321000000e-07 V_hig
+ 3.321010000e-07 V_hig
+ 3.322000000e-07 V_hig
+ 3.322010000e-07 V_hig
+ 3.323000000e-07 V_hig
+ 3.323010000e-07 V_hig
+ 3.324000000e-07 V_hig
+ 3.324010000e-07 V_hig
+ 3.325000000e-07 V_hig
+ 3.325010000e-07 V_hig
+ 3.326000000e-07 V_hig
+ 3.326010000e-07 V_hig
+ 3.327000000e-07 V_hig
+ 3.327010000e-07 V_hig
+ 3.328000000e-07 V_hig
+ 3.328010000e-07 V_hig
+ 3.329000000e-07 V_hig
+ 3.329010000e-07 V_low
+ 3.330000000e-07 V_low
+ 3.330010000e-07 V_low
+ 3.331000000e-07 V_low
+ 3.331010000e-07 V_low
+ 3.332000000e-07 V_low
+ 3.332010000e-07 V_low
+ 3.333000000e-07 V_low
+ 3.333010000e-07 V_low
+ 3.334000000e-07 V_low
+ 3.334010000e-07 V_low
+ 3.335000000e-07 V_low
+ 3.335010000e-07 V_low
+ 3.336000000e-07 V_low
+ 3.336010000e-07 V_low
+ 3.337000000e-07 V_low
+ 3.337010000e-07 V_low
+ 3.338000000e-07 V_low
+ 3.338010000e-07 V_low
+ 3.339000000e-07 V_low
+ 3.339010000e-07 V_low
+ 3.340000000e-07 V_low
+ 3.340010000e-07 V_low
+ 3.341000000e-07 V_low
+ 3.341010000e-07 V_low
+ 3.342000000e-07 V_low
+ 3.342010000e-07 V_low
+ 3.343000000e-07 V_low
+ 3.343010000e-07 V_low
+ 3.344000000e-07 V_low
+ 3.344010000e-07 V_low
+ 3.345000000e-07 V_low
+ 3.345010000e-07 V_low
+ 3.346000000e-07 V_low
+ 3.346010000e-07 V_low
+ 3.347000000e-07 V_low
+ 3.347010000e-07 V_low
+ 3.348000000e-07 V_low
+ 3.348010000e-07 V_low
+ 3.349000000e-07 V_low
+ 3.349010000e-07 V_low
+ 3.350000000e-07 V_low
+ 3.350010000e-07 V_low
+ 3.351000000e-07 V_low
+ 3.351010000e-07 V_low
+ 3.352000000e-07 V_low
+ 3.352010000e-07 V_low
+ 3.353000000e-07 V_low
+ 3.353010000e-07 V_low
+ 3.354000000e-07 V_low
+ 3.354010000e-07 V_low
+ 3.355000000e-07 V_low
+ 3.355010000e-07 V_low
+ 3.356000000e-07 V_low
+ 3.356010000e-07 V_low
+ 3.357000000e-07 V_low
+ 3.357010000e-07 V_low
+ 3.358000000e-07 V_low
+ 3.358010000e-07 V_low
+ 3.359000000e-07 V_low
+ 3.359010000e-07 V_hig
+ 3.360000000e-07 V_hig
+ 3.360010000e-07 V_hig
+ 3.361000000e-07 V_hig
+ 3.361010000e-07 V_hig
+ 3.362000000e-07 V_hig
+ 3.362010000e-07 V_hig
+ 3.363000000e-07 V_hig
+ 3.363010000e-07 V_hig
+ 3.364000000e-07 V_hig
+ 3.364010000e-07 V_hig
+ 3.365000000e-07 V_hig
+ 3.365010000e-07 V_hig
+ 3.366000000e-07 V_hig
+ 3.366010000e-07 V_hig
+ 3.367000000e-07 V_hig
+ 3.367010000e-07 V_hig
+ 3.368000000e-07 V_hig
+ 3.368010000e-07 V_hig
+ 3.369000000e-07 V_hig
+ 3.369010000e-07 V_low
+ 3.370000000e-07 V_low
+ 3.370010000e-07 V_low
+ 3.371000000e-07 V_low
+ 3.371010000e-07 V_low
+ 3.372000000e-07 V_low
+ 3.372010000e-07 V_low
+ 3.373000000e-07 V_low
+ 3.373010000e-07 V_low
+ 3.374000000e-07 V_low
+ 3.374010000e-07 V_low
+ 3.375000000e-07 V_low
+ 3.375010000e-07 V_low
+ 3.376000000e-07 V_low
+ 3.376010000e-07 V_low
+ 3.377000000e-07 V_low
+ 3.377010000e-07 V_low
+ 3.378000000e-07 V_low
+ 3.378010000e-07 V_low
+ 3.379000000e-07 V_low
+ 3.379010000e-07 V_low
+ 3.380000000e-07 V_low
+ 3.380010000e-07 V_low
+ 3.381000000e-07 V_low
+ 3.381010000e-07 V_low
+ 3.382000000e-07 V_low
+ 3.382010000e-07 V_low
+ 3.383000000e-07 V_low
+ 3.383010000e-07 V_low
+ 3.384000000e-07 V_low
+ 3.384010000e-07 V_low
+ 3.385000000e-07 V_low
+ 3.385010000e-07 V_low
+ 3.386000000e-07 V_low
+ 3.386010000e-07 V_low
+ 3.387000000e-07 V_low
+ 3.387010000e-07 V_low
+ 3.388000000e-07 V_low
+ 3.388010000e-07 V_low
+ 3.389000000e-07 V_low
+ 3.389010000e-07 V_low
+ 3.390000000e-07 V_low
+ 3.390010000e-07 V_low
+ 3.391000000e-07 V_low
+ 3.391010000e-07 V_low
+ 3.392000000e-07 V_low
+ 3.392010000e-07 V_low
+ 3.393000000e-07 V_low
+ 3.393010000e-07 V_low
+ 3.394000000e-07 V_low
+ 3.394010000e-07 V_low
+ 3.395000000e-07 V_low
+ 3.395010000e-07 V_low
+ 3.396000000e-07 V_low
+ 3.396010000e-07 V_low
+ 3.397000000e-07 V_low
+ 3.397010000e-07 V_low
+ 3.398000000e-07 V_low
+ 3.398010000e-07 V_low
+ 3.399000000e-07 V_low
+ 3.399010000e-07 V_low
+ 3.400000000e-07 V_low
+ 3.400010000e-07 V_low
+ 3.401000000e-07 V_low
+ 3.401010000e-07 V_low
+ 3.402000000e-07 V_low
+ 3.402010000e-07 V_low
+ 3.403000000e-07 V_low
+ 3.403010000e-07 V_low
+ 3.404000000e-07 V_low
+ 3.404010000e-07 V_low
+ 3.405000000e-07 V_low
+ 3.405010000e-07 V_low
+ 3.406000000e-07 V_low
+ 3.406010000e-07 V_low
+ 3.407000000e-07 V_low
+ 3.407010000e-07 V_low
+ 3.408000000e-07 V_low
+ 3.408010000e-07 V_low
+ 3.409000000e-07 V_low
+ 3.409010000e-07 V_hig
+ 3.410000000e-07 V_hig
+ 3.410010000e-07 V_hig
+ 3.411000000e-07 V_hig
+ 3.411010000e-07 V_hig
+ 3.412000000e-07 V_hig
+ 3.412010000e-07 V_hig
+ 3.413000000e-07 V_hig
+ 3.413010000e-07 V_hig
+ 3.414000000e-07 V_hig
+ 3.414010000e-07 V_hig
+ 3.415000000e-07 V_hig
+ 3.415010000e-07 V_hig
+ 3.416000000e-07 V_hig
+ 3.416010000e-07 V_hig
+ 3.417000000e-07 V_hig
+ 3.417010000e-07 V_hig
+ 3.418000000e-07 V_hig
+ 3.418010000e-07 V_hig
+ 3.419000000e-07 V_hig
+ 3.419010000e-07 V_hig
+ 3.420000000e-07 V_hig
+ 3.420010000e-07 V_hig
+ 3.421000000e-07 V_hig
+ 3.421010000e-07 V_hig
+ 3.422000000e-07 V_hig
+ 3.422010000e-07 V_hig
+ 3.423000000e-07 V_hig
+ 3.423010000e-07 V_hig
+ 3.424000000e-07 V_hig
+ 3.424010000e-07 V_hig
+ 3.425000000e-07 V_hig
+ 3.425010000e-07 V_hig
+ 3.426000000e-07 V_hig
+ 3.426010000e-07 V_hig
+ 3.427000000e-07 V_hig
+ 3.427010000e-07 V_hig
+ 3.428000000e-07 V_hig
+ 3.428010000e-07 V_hig
+ 3.429000000e-07 V_hig
+ 3.429010000e-07 V_hig
+ 3.430000000e-07 V_hig
+ 3.430010000e-07 V_hig
+ 3.431000000e-07 V_hig
+ 3.431010000e-07 V_hig
+ 3.432000000e-07 V_hig
+ 3.432010000e-07 V_hig
+ 3.433000000e-07 V_hig
+ 3.433010000e-07 V_hig
+ 3.434000000e-07 V_hig
+ 3.434010000e-07 V_hig
+ 3.435000000e-07 V_hig
+ 3.435010000e-07 V_hig
+ 3.436000000e-07 V_hig
+ 3.436010000e-07 V_hig
+ 3.437000000e-07 V_hig
+ 3.437010000e-07 V_hig
+ 3.438000000e-07 V_hig
+ 3.438010000e-07 V_hig
+ 3.439000000e-07 V_hig
+ 3.439010000e-07 V_low
+ 3.440000000e-07 V_low
+ 3.440010000e-07 V_low
+ 3.441000000e-07 V_low
+ 3.441010000e-07 V_low
+ 3.442000000e-07 V_low
+ 3.442010000e-07 V_low
+ 3.443000000e-07 V_low
+ 3.443010000e-07 V_low
+ 3.444000000e-07 V_low
+ 3.444010000e-07 V_low
+ 3.445000000e-07 V_low
+ 3.445010000e-07 V_low
+ 3.446000000e-07 V_low
+ 3.446010000e-07 V_low
+ 3.447000000e-07 V_low
+ 3.447010000e-07 V_low
+ 3.448000000e-07 V_low
+ 3.448010000e-07 V_low
+ 3.449000000e-07 V_low
+ 3.449010000e-07 V_hig
+ 3.450000000e-07 V_hig
+ 3.450010000e-07 V_hig
+ 3.451000000e-07 V_hig
+ 3.451010000e-07 V_hig
+ 3.452000000e-07 V_hig
+ 3.452010000e-07 V_hig
+ 3.453000000e-07 V_hig
+ 3.453010000e-07 V_hig
+ 3.454000000e-07 V_hig
+ 3.454010000e-07 V_hig
+ 3.455000000e-07 V_hig
+ 3.455010000e-07 V_hig
+ 3.456000000e-07 V_hig
+ 3.456010000e-07 V_hig
+ 3.457000000e-07 V_hig
+ 3.457010000e-07 V_hig
+ 3.458000000e-07 V_hig
+ 3.458010000e-07 V_hig
+ 3.459000000e-07 V_hig
+ 3.459010000e-07 V_low
+ 3.460000000e-07 V_low
+ 3.460010000e-07 V_low
+ 3.461000000e-07 V_low
+ 3.461010000e-07 V_low
+ 3.462000000e-07 V_low
+ 3.462010000e-07 V_low
+ 3.463000000e-07 V_low
+ 3.463010000e-07 V_low
+ 3.464000000e-07 V_low
+ 3.464010000e-07 V_low
+ 3.465000000e-07 V_low
+ 3.465010000e-07 V_low
+ 3.466000000e-07 V_low
+ 3.466010000e-07 V_low
+ 3.467000000e-07 V_low
+ 3.467010000e-07 V_low
+ 3.468000000e-07 V_low
+ 3.468010000e-07 V_low
+ 3.469000000e-07 V_low
+ 3.469010000e-07 V_low
+ 3.470000000e-07 V_low
+ 3.470010000e-07 V_low
+ 3.471000000e-07 V_low
+ 3.471010000e-07 V_low
+ 3.472000000e-07 V_low
+ 3.472010000e-07 V_low
+ 3.473000000e-07 V_low
+ 3.473010000e-07 V_low
+ 3.474000000e-07 V_low
+ 3.474010000e-07 V_low
+ 3.475000000e-07 V_low
+ 3.475010000e-07 V_low
+ 3.476000000e-07 V_low
+ 3.476010000e-07 V_low
+ 3.477000000e-07 V_low
+ 3.477010000e-07 V_low
+ 3.478000000e-07 V_low
+ 3.478010000e-07 V_low
+ 3.479000000e-07 V_low
+ 3.479010000e-07 V_low
+ 3.480000000e-07 V_low
+ 3.480010000e-07 V_low
+ 3.481000000e-07 V_low
+ 3.481010000e-07 V_low
+ 3.482000000e-07 V_low
+ 3.482010000e-07 V_low
+ 3.483000000e-07 V_low
+ 3.483010000e-07 V_low
+ 3.484000000e-07 V_low
+ 3.484010000e-07 V_low
+ 3.485000000e-07 V_low
+ 3.485010000e-07 V_low
+ 3.486000000e-07 V_low
+ 3.486010000e-07 V_low
+ 3.487000000e-07 V_low
+ 3.487010000e-07 V_low
+ 3.488000000e-07 V_low
+ 3.488010000e-07 V_low
+ 3.489000000e-07 V_low
+ 3.489010000e-07 V_low
+ 3.490000000e-07 V_low
+ 3.490010000e-07 V_low
+ 3.491000000e-07 V_low
+ 3.491010000e-07 V_low
+ 3.492000000e-07 V_low
+ 3.492010000e-07 V_low
+ 3.493000000e-07 V_low
+ 3.493010000e-07 V_low
+ 3.494000000e-07 V_low
+ 3.494010000e-07 V_low
+ 3.495000000e-07 V_low
+ 3.495010000e-07 V_low
+ 3.496000000e-07 V_low
+ 3.496010000e-07 V_low
+ 3.497000000e-07 V_low
+ 3.497010000e-07 V_low
+ 3.498000000e-07 V_low
+ 3.498010000e-07 V_low
+ 3.499000000e-07 V_low
+ 3.499010000e-07 V_hig
+ 3.500000000e-07 V_hig
+ 3.500010000e-07 V_hig
+ 3.501000000e-07 V_hig
+ 3.501010000e-07 V_hig
+ 3.502000000e-07 V_hig
+ 3.502010000e-07 V_hig
+ 3.503000000e-07 V_hig
+ 3.503010000e-07 V_hig
+ 3.504000000e-07 V_hig
+ 3.504010000e-07 V_hig
+ 3.505000000e-07 V_hig
+ 3.505010000e-07 V_hig
+ 3.506000000e-07 V_hig
+ 3.506010000e-07 V_hig
+ 3.507000000e-07 V_hig
+ 3.507010000e-07 V_hig
+ 3.508000000e-07 V_hig
+ 3.508010000e-07 V_hig
+ 3.509000000e-07 V_hig
+ 3.509010000e-07 V_low
+ 3.510000000e-07 V_low
+ 3.510010000e-07 V_low
+ 3.511000000e-07 V_low
+ 3.511010000e-07 V_low
+ 3.512000000e-07 V_low
+ 3.512010000e-07 V_low
+ 3.513000000e-07 V_low
+ 3.513010000e-07 V_low
+ 3.514000000e-07 V_low
+ 3.514010000e-07 V_low
+ 3.515000000e-07 V_low
+ 3.515010000e-07 V_low
+ 3.516000000e-07 V_low
+ 3.516010000e-07 V_low
+ 3.517000000e-07 V_low
+ 3.517010000e-07 V_low
+ 3.518000000e-07 V_low
+ 3.518010000e-07 V_low
+ 3.519000000e-07 V_low
+ 3.519010000e-07 V_hig
+ 3.520000000e-07 V_hig
+ 3.520010000e-07 V_hig
+ 3.521000000e-07 V_hig
+ 3.521010000e-07 V_hig
+ 3.522000000e-07 V_hig
+ 3.522010000e-07 V_hig
+ 3.523000000e-07 V_hig
+ 3.523010000e-07 V_hig
+ 3.524000000e-07 V_hig
+ 3.524010000e-07 V_hig
+ 3.525000000e-07 V_hig
+ 3.525010000e-07 V_hig
+ 3.526000000e-07 V_hig
+ 3.526010000e-07 V_hig
+ 3.527000000e-07 V_hig
+ 3.527010000e-07 V_hig
+ 3.528000000e-07 V_hig
+ 3.528010000e-07 V_hig
+ 3.529000000e-07 V_hig
+ 3.529010000e-07 V_hig
+ 3.530000000e-07 V_hig
+ 3.530010000e-07 V_hig
+ 3.531000000e-07 V_hig
+ 3.531010000e-07 V_hig
+ 3.532000000e-07 V_hig
+ 3.532010000e-07 V_hig
+ 3.533000000e-07 V_hig
+ 3.533010000e-07 V_hig
+ 3.534000000e-07 V_hig
+ 3.534010000e-07 V_hig
+ 3.535000000e-07 V_hig
+ 3.535010000e-07 V_hig
+ 3.536000000e-07 V_hig
+ 3.536010000e-07 V_hig
+ 3.537000000e-07 V_hig
+ 3.537010000e-07 V_hig
+ 3.538000000e-07 V_hig
+ 3.538010000e-07 V_hig
+ 3.539000000e-07 V_hig
+ 3.539010000e-07 V_hig
+ 3.540000000e-07 V_hig
+ 3.540010000e-07 V_hig
+ 3.541000000e-07 V_hig
+ 3.541010000e-07 V_hig
+ 3.542000000e-07 V_hig
+ 3.542010000e-07 V_hig
+ 3.543000000e-07 V_hig
+ 3.543010000e-07 V_hig
+ 3.544000000e-07 V_hig
+ 3.544010000e-07 V_hig
+ 3.545000000e-07 V_hig
+ 3.545010000e-07 V_hig
+ 3.546000000e-07 V_hig
+ 3.546010000e-07 V_hig
+ 3.547000000e-07 V_hig
+ 3.547010000e-07 V_hig
+ 3.548000000e-07 V_hig
+ 3.548010000e-07 V_hig
+ 3.549000000e-07 V_hig
+ 3.549010000e-07 V_low
+ 3.550000000e-07 V_low
+ 3.550010000e-07 V_low
+ 3.551000000e-07 V_low
+ 3.551010000e-07 V_low
+ 3.552000000e-07 V_low
+ 3.552010000e-07 V_low
+ 3.553000000e-07 V_low
+ 3.553010000e-07 V_low
+ 3.554000000e-07 V_low
+ 3.554010000e-07 V_low
+ 3.555000000e-07 V_low
+ 3.555010000e-07 V_low
+ 3.556000000e-07 V_low
+ 3.556010000e-07 V_low
+ 3.557000000e-07 V_low
+ 3.557010000e-07 V_low
+ 3.558000000e-07 V_low
+ 3.558010000e-07 V_low
+ 3.559000000e-07 V_low
+ 3.559010000e-07 V_low
+ 3.560000000e-07 V_low
+ 3.560010000e-07 V_low
+ 3.561000000e-07 V_low
+ 3.561010000e-07 V_low
+ 3.562000000e-07 V_low
+ 3.562010000e-07 V_low
+ 3.563000000e-07 V_low
+ 3.563010000e-07 V_low
+ 3.564000000e-07 V_low
+ 3.564010000e-07 V_low
+ 3.565000000e-07 V_low
+ 3.565010000e-07 V_low
+ 3.566000000e-07 V_low
+ 3.566010000e-07 V_low
+ 3.567000000e-07 V_low
+ 3.567010000e-07 V_low
+ 3.568000000e-07 V_low
+ 3.568010000e-07 V_low
+ 3.569000000e-07 V_low
+ 3.569010000e-07 V_low
+ 3.570000000e-07 V_low
+ 3.570010000e-07 V_low
+ 3.571000000e-07 V_low
+ 3.571010000e-07 V_low
+ 3.572000000e-07 V_low
+ 3.572010000e-07 V_low
+ 3.573000000e-07 V_low
+ 3.573010000e-07 V_low
+ 3.574000000e-07 V_low
+ 3.574010000e-07 V_low
+ 3.575000000e-07 V_low
+ 3.575010000e-07 V_low
+ 3.576000000e-07 V_low
+ 3.576010000e-07 V_low
+ 3.577000000e-07 V_low
+ 3.577010000e-07 V_low
+ 3.578000000e-07 V_low
+ 3.578010000e-07 V_low
+ 3.579000000e-07 V_low
+ 3.579010000e-07 V_hig
+ 3.580000000e-07 V_hig
+ 3.580010000e-07 V_hig
+ 3.581000000e-07 V_hig
+ 3.581010000e-07 V_hig
+ 3.582000000e-07 V_hig
+ 3.582010000e-07 V_hig
+ 3.583000000e-07 V_hig
+ 3.583010000e-07 V_hig
+ 3.584000000e-07 V_hig
+ 3.584010000e-07 V_hig
+ 3.585000000e-07 V_hig
+ 3.585010000e-07 V_hig
+ 3.586000000e-07 V_hig
+ 3.586010000e-07 V_hig
+ 3.587000000e-07 V_hig
+ 3.587010000e-07 V_hig
+ 3.588000000e-07 V_hig
+ 3.588010000e-07 V_hig
+ 3.589000000e-07 V_hig
+ 3.589010000e-07 V_low
+ 3.590000000e-07 V_low
+ 3.590010000e-07 V_low
+ 3.591000000e-07 V_low
+ 3.591010000e-07 V_low
+ 3.592000000e-07 V_low
+ 3.592010000e-07 V_low
+ 3.593000000e-07 V_low
+ 3.593010000e-07 V_low
+ 3.594000000e-07 V_low
+ 3.594010000e-07 V_low
+ 3.595000000e-07 V_low
+ 3.595010000e-07 V_low
+ 3.596000000e-07 V_low
+ 3.596010000e-07 V_low
+ 3.597000000e-07 V_low
+ 3.597010000e-07 V_low
+ 3.598000000e-07 V_low
+ 3.598010000e-07 V_low
+ 3.599000000e-07 V_low
+ 3.599010000e-07 V_hig
+ 3.600000000e-07 V_hig
+ 3.600010000e-07 V_hig
+ 3.601000000e-07 V_hig
+ 3.601010000e-07 V_hig
+ 3.602000000e-07 V_hig
+ 3.602010000e-07 V_hig
+ 3.603000000e-07 V_hig
+ 3.603010000e-07 V_hig
+ 3.604000000e-07 V_hig
+ 3.604010000e-07 V_hig
+ 3.605000000e-07 V_hig
+ 3.605010000e-07 V_hig
+ 3.606000000e-07 V_hig
+ 3.606010000e-07 V_hig
+ 3.607000000e-07 V_hig
+ 3.607010000e-07 V_hig
+ 3.608000000e-07 V_hig
+ 3.608010000e-07 V_hig
+ 3.609000000e-07 V_hig
+ 3.609010000e-07 V_low
+ 3.610000000e-07 V_low
+ 3.610010000e-07 V_low
+ 3.611000000e-07 V_low
+ 3.611010000e-07 V_low
+ 3.612000000e-07 V_low
+ 3.612010000e-07 V_low
+ 3.613000000e-07 V_low
+ 3.613010000e-07 V_low
+ 3.614000000e-07 V_low
+ 3.614010000e-07 V_low
+ 3.615000000e-07 V_low
+ 3.615010000e-07 V_low
+ 3.616000000e-07 V_low
+ 3.616010000e-07 V_low
+ 3.617000000e-07 V_low
+ 3.617010000e-07 V_low
+ 3.618000000e-07 V_low
+ 3.618010000e-07 V_low
+ 3.619000000e-07 V_low
+ 3.619010000e-07 V_hig
+ 3.620000000e-07 V_hig
+ 3.620010000e-07 V_hig
+ 3.621000000e-07 V_hig
+ 3.621010000e-07 V_hig
+ 3.622000000e-07 V_hig
+ 3.622010000e-07 V_hig
+ 3.623000000e-07 V_hig
+ 3.623010000e-07 V_hig
+ 3.624000000e-07 V_hig
+ 3.624010000e-07 V_hig
+ 3.625000000e-07 V_hig
+ 3.625010000e-07 V_hig
+ 3.626000000e-07 V_hig
+ 3.626010000e-07 V_hig
+ 3.627000000e-07 V_hig
+ 3.627010000e-07 V_hig
+ 3.628000000e-07 V_hig
+ 3.628010000e-07 V_hig
+ 3.629000000e-07 V_hig
+ 3.629010000e-07 V_low
+ 3.630000000e-07 V_low
+ 3.630010000e-07 V_low
+ 3.631000000e-07 V_low
+ 3.631010000e-07 V_low
+ 3.632000000e-07 V_low
+ 3.632010000e-07 V_low
+ 3.633000000e-07 V_low
+ 3.633010000e-07 V_low
+ 3.634000000e-07 V_low
+ 3.634010000e-07 V_low
+ 3.635000000e-07 V_low
+ 3.635010000e-07 V_low
+ 3.636000000e-07 V_low
+ 3.636010000e-07 V_low
+ 3.637000000e-07 V_low
+ 3.637010000e-07 V_low
+ 3.638000000e-07 V_low
+ 3.638010000e-07 V_low
+ 3.639000000e-07 V_low
+ 3.639010000e-07 V_low
+ 3.640000000e-07 V_low
+ 3.640010000e-07 V_low
+ 3.641000000e-07 V_low
+ 3.641010000e-07 V_low
+ 3.642000000e-07 V_low
+ 3.642010000e-07 V_low
+ 3.643000000e-07 V_low
+ 3.643010000e-07 V_low
+ 3.644000000e-07 V_low
+ 3.644010000e-07 V_low
+ 3.645000000e-07 V_low
+ 3.645010000e-07 V_low
+ 3.646000000e-07 V_low
+ 3.646010000e-07 V_low
+ 3.647000000e-07 V_low
+ 3.647010000e-07 V_low
+ 3.648000000e-07 V_low
+ 3.648010000e-07 V_low
+ 3.649000000e-07 V_low
+ 3.649010000e-07 V_hig
+ 3.650000000e-07 V_hig
+ 3.650010000e-07 V_hig
+ 3.651000000e-07 V_hig
+ 3.651010000e-07 V_hig
+ 3.652000000e-07 V_hig
+ 3.652010000e-07 V_hig
+ 3.653000000e-07 V_hig
+ 3.653010000e-07 V_hig
+ 3.654000000e-07 V_hig
+ 3.654010000e-07 V_hig
+ 3.655000000e-07 V_hig
+ 3.655010000e-07 V_hig
+ 3.656000000e-07 V_hig
+ 3.656010000e-07 V_hig
+ 3.657000000e-07 V_hig
+ 3.657010000e-07 V_hig
+ 3.658000000e-07 V_hig
+ 3.658010000e-07 V_hig
+ 3.659000000e-07 V_hig
+ 3.659010000e-07 V_low
+ 3.660000000e-07 V_low
+ 3.660010000e-07 V_low
+ 3.661000000e-07 V_low
+ 3.661010000e-07 V_low
+ 3.662000000e-07 V_low
+ 3.662010000e-07 V_low
+ 3.663000000e-07 V_low
+ 3.663010000e-07 V_low
+ 3.664000000e-07 V_low
+ 3.664010000e-07 V_low
+ 3.665000000e-07 V_low
+ 3.665010000e-07 V_low
+ 3.666000000e-07 V_low
+ 3.666010000e-07 V_low
+ 3.667000000e-07 V_low
+ 3.667010000e-07 V_low
+ 3.668000000e-07 V_low
+ 3.668010000e-07 V_low
+ 3.669000000e-07 V_low
+ 3.669010000e-07 V_low
+ 3.670000000e-07 V_low
+ 3.670010000e-07 V_low
+ 3.671000000e-07 V_low
+ 3.671010000e-07 V_low
+ 3.672000000e-07 V_low
+ 3.672010000e-07 V_low
+ 3.673000000e-07 V_low
+ 3.673010000e-07 V_low
+ 3.674000000e-07 V_low
+ 3.674010000e-07 V_low
+ 3.675000000e-07 V_low
+ 3.675010000e-07 V_low
+ 3.676000000e-07 V_low
+ 3.676010000e-07 V_low
+ 3.677000000e-07 V_low
+ 3.677010000e-07 V_low
+ 3.678000000e-07 V_low
+ 3.678010000e-07 V_low
+ 3.679000000e-07 V_low
+ 3.679010000e-07 V_hig
+ 3.680000000e-07 V_hig
+ 3.680010000e-07 V_hig
+ 3.681000000e-07 V_hig
+ 3.681010000e-07 V_hig
+ 3.682000000e-07 V_hig
+ 3.682010000e-07 V_hig
+ 3.683000000e-07 V_hig
+ 3.683010000e-07 V_hig
+ 3.684000000e-07 V_hig
+ 3.684010000e-07 V_hig
+ 3.685000000e-07 V_hig
+ 3.685010000e-07 V_hig
+ 3.686000000e-07 V_hig
+ 3.686010000e-07 V_hig
+ 3.687000000e-07 V_hig
+ 3.687010000e-07 V_hig
+ 3.688000000e-07 V_hig
+ 3.688010000e-07 V_hig
+ 3.689000000e-07 V_hig
+ 3.689010000e-07 V_hig
+ 3.690000000e-07 V_hig
+ 3.690010000e-07 V_hig
+ 3.691000000e-07 V_hig
+ 3.691010000e-07 V_hig
+ 3.692000000e-07 V_hig
+ 3.692010000e-07 V_hig
+ 3.693000000e-07 V_hig
+ 3.693010000e-07 V_hig
+ 3.694000000e-07 V_hig
+ 3.694010000e-07 V_hig
+ 3.695000000e-07 V_hig
+ 3.695010000e-07 V_hig
+ 3.696000000e-07 V_hig
+ 3.696010000e-07 V_hig
+ 3.697000000e-07 V_hig
+ 3.697010000e-07 V_hig
+ 3.698000000e-07 V_hig
+ 3.698010000e-07 V_hig
+ 3.699000000e-07 V_hig
+ 3.699010000e-07 V_low
+ 3.700000000e-07 V_low
+ 3.700010000e-07 V_low
+ 3.701000000e-07 V_low
+ 3.701010000e-07 V_low
+ 3.702000000e-07 V_low
+ 3.702010000e-07 V_low
+ 3.703000000e-07 V_low
+ 3.703010000e-07 V_low
+ 3.704000000e-07 V_low
+ 3.704010000e-07 V_low
+ 3.705000000e-07 V_low
+ 3.705010000e-07 V_low
+ 3.706000000e-07 V_low
+ 3.706010000e-07 V_low
+ 3.707000000e-07 V_low
+ 3.707010000e-07 V_low
+ 3.708000000e-07 V_low
+ 3.708010000e-07 V_low
+ 3.709000000e-07 V_low
+ 3.709010000e-07 V_hig
+ 3.710000000e-07 V_hig
+ 3.710010000e-07 V_hig
+ 3.711000000e-07 V_hig
+ 3.711010000e-07 V_hig
+ 3.712000000e-07 V_hig
+ 3.712010000e-07 V_hig
+ 3.713000000e-07 V_hig
+ 3.713010000e-07 V_hig
+ 3.714000000e-07 V_hig
+ 3.714010000e-07 V_hig
+ 3.715000000e-07 V_hig
+ 3.715010000e-07 V_hig
+ 3.716000000e-07 V_hig
+ 3.716010000e-07 V_hig
+ 3.717000000e-07 V_hig
+ 3.717010000e-07 V_hig
+ 3.718000000e-07 V_hig
+ 3.718010000e-07 V_hig
+ 3.719000000e-07 V_hig
+ 3.719010000e-07 V_low
+ 3.720000000e-07 V_low
+ 3.720010000e-07 V_low
+ 3.721000000e-07 V_low
+ 3.721010000e-07 V_low
+ 3.722000000e-07 V_low
+ 3.722010000e-07 V_low
+ 3.723000000e-07 V_low
+ 3.723010000e-07 V_low
+ 3.724000000e-07 V_low
+ 3.724010000e-07 V_low
+ 3.725000000e-07 V_low
+ 3.725010000e-07 V_low
+ 3.726000000e-07 V_low
+ 3.726010000e-07 V_low
+ 3.727000000e-07 V_low
+ 3.727010000e-07 V_low
+ 3.728000000e-07 V_low
+ 3.728010000e-07 V_low
+ 3.729000000e-07 V_low
+ 3.729010000e-07 V_low
+ 3.730000000e-07 V_low
+ 3.730010000e-07 V_low
+ 3.731000000e-07 V_low
+ 3.731010000e-07 V_low
+ 3.732000000e-07 V_low
+ 3.732010000e-07 V_low
+ 3.733000000e-07 V_low
+ 3.733010000e-07 V_low
+ 3.734000000e-07 V_low
+ 3.734010000e-07 V_low
+ 3.735000000e-07 V_low
+ 3.735010000e-07 V_low
+ 3.736000000e-07 V_low
+ 3.736010000e-07 V_low
+ 3.737000000e-07 V_low
+ 3.737010000e-07 V_low
+ 3.738000000e-07 V_low
+ 3.738010000e-07 V_low
+ 3.739000000e-07 V_low
+ 3.739010000e-07 V_low
+ 3.740000000e-07 V_low
+ 3.740010000e-07 V_low
+ 3.741000000e-07 V_low
+ 3.741010000e-07 V_low
+ 3.742000000e-07 V_low
+ 3.742010000e-07 V_low
+ 3.743000000e-07 V_low
+ 3.743010000e-07 V_low
+ 3.744000000e-07 V_low
+ 3.744010000e-07 V_low
+ 3.745000000e-07 V_low
+ 3.745010000e-07 V_low
+ 3.746000000e-07 V_low
+ 3.746010000e-07 V_low
+ 3.747000000e-07 V_low
+ 3.747010000e-07 V_low
+ 3.748000000e-07 V_low
+ 3.748010000e-07 V_low
+ 3.749000000e-07 V_low
+ 3.749010000e-07 V_low
+ 3.750000000e-07 V_low
+ 3.750010000e-07 V_low
+ 3.751000000e-07 V_low
+ 3.751010000e-07 V_low
+ 3.752000000e-07 V_low
+ 3.752010000e-07 V_low
+ 3.753000000e-07 V_low
+ 3.753010000e-07 V_low
+ 3.754000000e-07 V_low
+ 3.754010000e-07 V_low
+ 3.755000000e-07 V_low
+ 3.755010000e-07 V_low
+ 3.756000000e-07 V_low
+ 3.756010000e-07 V_low
+ 3.757000000e-07 V_low
+ 3.757010000e-07 V_low
+ 3.758000000e-07 V_low
+ 3.758010000e-07 V_low
+ 3.759000000e-07 V_low
+ 3.759010000e-07 V_hig
+ 3.760000000e-07 V_hig
+ 3.760010000e-07 V_hig
+ 3.761000000e-07 V_hig
+ 3.761010000e-07 V_hig
+ 3.762000000e-07 V_hig
+ 3.762010000e-07 V_hig
+ 3.763000000e-07 V_hig
+ 3.763010000e-07 V_hig
+ 3.764000000e-07 V_hig
+ 3.764010000e-07 V_hig
+ 3.765000000e-07 V_hig
+ 3.765010000e-07 V_hig
+ 3.766000000e-07 V_hig
+ 3.766010000e-07 V_hig
+ 3.767000000e-07 V_hig
+ 3.767010000e-07 V_hig
+ 3.768000000e-07 V_hig
+ 3.768010000e-07 V_hig
+ 3.769000000e-07 V_hig
+ 3.769010000e-07 V_low
+ 3.770000000e-07 V_low
+ 3.770010000e-07 V_low
+ 3.771000000e-07 V_low
+ 3.771010000e-07 V_low
+ 3.772000000e-07 V_low
+ 3.772010000e-07 V_low
+ 3.773000000e-07 V_low
+ 3.773010000e-07 V_low
+ 3.774000000e-07 V_low
+ 3.774010000e-07 V_low
+ 3.775000000e-07 V_low
+ 3.775010000e-07 V_low
+ 3.776000000e-07 V_low
+ 3.776010000e-07 V_low
+ 3.777000000e-07 V_low
+ 3.777010000e-07 V_low
+ 3.778000000e-07 V_low
+ 3.778010000e-07 V_low
+ 3.779000000e-07 V_low
+ 3.779010000e-07 V_hig
+ 3.780000000e-07 V_hig
+ 3.780010000e-07 V_hig
+ 3.781000000e-07 V_hig
+ 3.781010000e-07 V_hig
+ 3.782000000e-07 V_hig
+ 3.782010000e-07 V_hig
+ 3.783000000e-07 V_hig
+ 3.783010000e-07 V_hig
+ 3.784000000e-07 V_hig
+ 3.784010000e-07 V_hig
+ 3.785000000e-07 V_hig
+ 3.785010000e-07 V_hig
+ 3.786000000e-07 V_hig
+ 3.786010000e-07 V_hig
+ 3.787000000e-07 V_hig
+ 3.787010000e-07 V_hig
+ 3.788000000e-07 V_hig
+ 3.788010000e-07 V_hig
+ 3.789000000e-07 V_hig
+ 3.789010000e-07 V_hig
+ 3.790000000e-07 V_hig
+ 3.790010000e-07 V_hig
+ 3.791000000e-07 V_hig
+ 3.791010000e-07 V_hig
+ 3.792000000e-07 V_hig
+ 3.792010000e-07 V_hig
+ 3.793000000e-07 V_hig
+ 3.793010000e-07 V_hig
+ 3.794000000e-07 V_hig
+ 3.794010000e-07 V_hig
+ 3.795000000e-07 V_hig
+ 3.795010000e-07 V_hig
+ 3.796000000e-07 V_hig
+ 3.796010000e-07 V_hig
+ 3.797000000e-07 V_hig
+ 3.797010000e-07 V_hig
+ 3.798000000e-07 V_hig
+ 3.798010000e-07 V_hig
+ 3.799000000e-07 V_hig
+ 3.799010000e-07 V_low
+ 3.800000000e-07 V_low
+ 3.800010000e-07 V_low
+ 3.801000000e-07 V_low
+ 3.801010000e-07 V_low
+ 3.802000000e-07 V_low
+ 3.802010000e-07 V_low
+ 3.803000000e-07 V_low
+ 3.803010000e-07 V_low
+ 3.804000000e-07 V_low
+ 3.804010000e-07 V_low
+ 3.805000000e-07 V_low
+ 3.805010000e-07 V_low
+ 3.806000000e-07 V_low
+ 3.806010000e-07 V_low
+ 3.807000000e-07 V_low
+ 3.807010000e-07 V_low
+ 3.808000000e-07 V_low
+ 3.808010000e-07 V_low
+ 3.809000000e-07 V_low
+ 3.809010000e-07 V_hig
+ 3.810000000e-07 V_hig
+ 3.810010000e-07 V_hig
+ 3.811000000e-07 V_hig
+ 3.811010000e-07 V_hig
+ 3.812000000e-07 V_hig
+ 3.812010000e-07 V_hig
+ 3.813000000e-07 V_hig
+ 3.813010000e-07 V_hig
+ 3.814000000e-07 V_hig
+ 3.814010000e-07 V_hig
+ 3.815000000e-07 V_hig
+ 3.815010000e-07 V_hig
+ 3.816000000e-07 V_hig
+ 3.816010000e-07 V_hig
+ 3.817000000e-07 V_hig
+ 3.817010000e-07 V_hig
+ 3.818000000e-07 V_hig
+ 3.818010000e-07 V_hig
+ 3.819000000e-07 V_hig
+ 3.819010000e-07 V_hig
+ 3.820000000e-07 V_hig
+ 3.820010000e-07 V_hig
+ 3.821000000e-07 V_hig
+ 3.821010000e-07 V_hig
+ 3.822000000e-07 V_hig
+ 3.822010000e-07 V_hig
+ 3.823000000e-07 V_hig
+ 3.823010000e-07 V_hig
+ 3.824000000e-07 V_hig
+ 3.824010000e-07 V_hig
+ 3.825000000e-07 V_hig
+ 3.825010000e-07 V_hig
+ 3.826000000e-07 V_hig
+ 3.826010000e-07 V_hig
+ 3.827000000e-07 V_hig
+ 3.827010000e-07 V_hig
+ 3.828000000e-07 V_hig
+ 3.828010000e-07 V_hig
+ 3.829000000e-07 V_hig
+ 3.829010000e-07 V_low
+ 3.830000000e-07 V_low
+ 3.830010000e-07 V_low
+ 3.831000000e-07 V_low
+ 3.831010000e-07 V_low
+ 3.832000000e-07 V_low
+ 3.832010000e-07 V_low
+ 3.833000000e-07 V_low
+ 3.833010000e-07 V_low
+ 3.834000000e-07 V_low
+ 3.834010000e-07 V_low
+ 3.835000000e-07 V_low
+ 3.835010000e-07 V_low
+ 3.836000000e-07 V_low
+ 3.836010000e-07 V_low
+ 3.837000000e-07 V_low
+ 3.837010000e-07 V_low
+ 3.838000000e-07 V_low
+ 3.838010000e-07 V_low
+ 3.839000000e-07 V_low
+ 3.839010000e-07 V_hig
+ 3.840000000e-07 V_hig
+ 3.840010000e-07 V_hig
+ 3.841000000e-07 V_hig
+ 3.841010000e-07 V_hig
+ 3.842000000e-07 V_hig
+ 3.842010000e-07 V_hig
+ 3.843000000e-07 V_hig
+ 3.843010000e-07 V_hig
+ 3.844000000e-07 V_hig
+ 3.844010000e-07 V_hig
+ 3.845000000e-07 V_hig
+ 3.845010000e-07 V_hig
+ 3.846000000e-07 V_hig
+ 3.846010000e-07 V_hig
+ 3.847000000e-07 V_hig
+ 3.847010000e-07 V_hig
+ 3.848000000e-07 V_hig
+ 3.848010000e-07 V_hig
+ 3.849000000e-07 V_hig
+ 3.849010000e-07 V_low
+ 3.850000000e-07 V_low
+ 3.850010000e-07 V_low
+ 3.851000000e-07 V_low
+ 3.851010000e-07 V_low
+ 3.852000000e-07 V_low
+ 3.852010000e-07 V_low
+ 3.853000000e-07 V_low
+ 3.853010000e-07 V_low
+ 3.854000000e-07 V_low
+ 3.854010000e-07 V_low
+ 3.855000000e-07 V_low
+ 3.855010000e-07 V_low
+ 3.856000000e-07 V_low
+ 3.856010000e-07 V_low
+ 3.857000000e-07 V_low
+ 3.857010000e-07 V_low
+ 3.858000000e-07 V_low
+ 3.858010000e-07 V_low
+ 3.859000000e-07 V_low
+ 3.859010000e-07 V_hig
+ 3.860000000e-07 V_hig
+ 3.860010000e-07 V_hig
+ 3.861000000e-07 V_hig
+ 3.861010000e-07 V_hig
+ 3.862000000e-07 V_hig
+ 3.862010000e-07 V_hig
+ 3.863000000e-07 V_hig
+ 3.863010000e-07 V_hig
+ 3.864000000e-07 V_hig
+ 3.864010000e-07 V_hig
+ 3.865000000e-07 V_hig
+ 3.865010000e-07 V_hig
+ 3.866000000e-07 V_hig
+ 3.866010000e-07 V_hig
+ 3.867000000e-07 V_hig
+ 3.867010000e-07 V_hig
+ 3.868000000e-07 V_hig
+ 3.868010000e-07 V_hig
+ 3.869000000e-07 V_hig
+ 3.869010000e-07 V_low
+ 3.870000000e-07 V_low
+ 3.870010000e-07 V_low
+ 3.871000000e-07 V_low
+ 3.871010000e-07 V_low
+ 3.872000000e-07 V_low
+ 3.872010000e-07 V_low
+ 3.873000000e-07 V_low
+ 3.873010000e-07 V_low
+ 3.874000000e-07 V_low
+ 3.874010000e-07 V_low
+ 3.875000000e-07 V_low
+ 3.875010000e-07 V_low
+ 3.876000000e-07 V_low
+ 3.876010000e-07 V_low
+ 3.877000000e-07 V_low
+ 3.877010000e-07 V_low
+ 3.878000000e-07 V_low
+ 3.878010000e-07 V_low
+ 3.879000000e-07 V_low
+ 3.879010000e-07 V_low
+ 3.880000000e-07 V_low
+ 3.880010000e-07 V_low
+ 3.881000000e-07 V_low
+ 3.881010000e-07 V_low
+ 3.882000000e-07 V_low
+ 3.882010000e-07 V_low
+ 3.883000000e-07 V_low
+ 3.883010000e-07 V_low
+ 3.884000000e-07 V_low
+ 3.884010000e-07 V_low
+ 3.885000000e-07 V_low
+ 3.885010000e-07 V_low
+ 3.886000000e-07 V_low
+ 3.886010000e-07 V_low
+ 3.887000000e-07 V_low
+ 3.887010000e-07 V_low
+ 3.888000000e-07 V_low
+ 3.888010000e-07 V_low
+ 3.889000000e-07 V_low
+ 3.889010000e-07 V_hig
+ 3.890000000e-07 V_hig
+ 3.890010000e-07 V_hig
+ 3.891000000e-07 V_hig
+ 3.891010000e-07 V_hig
+ 3.892000000e-07 V_hig
+ 3.892010000e-07 V_hig
+ 3.893000000e-07 V_hig
+ 3.893010000e-07 V_hig
+ 3.894000000e-07 V_hig
+ 3.894010000e-07 V_hig
+ 3.895000000e-07 V_hig
+ 3.895010000e-07 V_hig
+ 3.896000000e-07 V_hig
+ 3.896010000e-07 V_hig
+ 3.897000000e-07 V_hig
+ 3.897010000e-07 V_hig
+ 3.898000000e-07 V_hig
+ 3.898010000e-07 V_hig
+ 3.899000000e-07 V_hig
+ 3.899010000e-07 V_hig
+ 3.900000000e-07 V_hig
+ 3.900010000e-07 V_hig
+ 3.901000000e-07 V_hig
+ 3.901010000e-07 V_hig
+ 3.902000000e-07 V_hig
+ 3.902010000e-07 V_hig
+ 3.903000000e-07 V_hig
+ 3.903010000e-07 V_hig
+ 3.904000000e-07 V_hig
+ 3.904010000e-07 V_hig
+ 3.905000000e-07 V_hig
+ 3.905010000e-07 V_hig
+ 3.906000000e-07 V_hig
+ 3.906010000e-07 V_hig
+ 3.907000000e-07 V_hig
+ 3.907010000e-07 V_hig
+ 3.908000000e-07 V_hig
+ 3.908010000e-07 V_hig
+ 3.909000000e-07 V_hig
+ 3.909010000e-07 V_hig
+ 3.910000000e-07 V_hig
+ 3.910010000e-07 V_hig
+ 3.911000000e-07 V_hig
+ 3.911010000e-07 V_hig
+ 3.912000000e-07 V_hig
+ 3.912010000e-07 V_hig
+ 3.913000000e-07 V_hig
+ 3.913010000e-07 V_hig
+ 3.914000000e-07 V_hig
+ 3.914010000e-07 V_hig
+ 3.915000000e-07 V_hig
+ 3.915010000e-07 V_hig
+ 3.916000000e-07 V_hig
+ 3.916010000e-07 V_hig
+ 3.917000000e-07 V_hig
+ 3.917010000e-07 V_hig
+ 3.918000000e-07 V_hig
+ 3.918010000e-07 V_hig
+ 3.919000000e-07 V_hig
+ 3.919010000e-07 V_hig
+ 3.920000000e-07 V_hig
+ 3.920010000e-07 V_hig
+ 3.921000000e-07 V_hig
+ 3.921010000e-07 V_hig
+ 3.922000000e-07 V_hig
+ 3.922010000e-07 V_hig
+ 3.923000000e-07 V_hig
+ 3.923010000e-07 V_hig
+ 3.924000000e-07 V_hig
+ 3.924010000e-07 V_hig
+ 3.925000000e-07 V_hig
+ 3.925010000e-07 V_hig
+ 3.926000000e-07 V_hig
+ 3.926010000e-07 V_hig
+ 3.927000000e-07 V_hig
+ 3.927010000e-07 V_hig
+ 3.928000000e-07 V_hig
+ 3.928010000e-07 V_hig
+ 3.929000000e-07 V_hig
+ 3.929010000e-07 V_low
+ 3.930000000e-07 V_low
+ 3.930010000e-07 V_low
+ 3.931000000e-07 V_low
+ 3.931010000e-07 V_low
+ 3.932000000e-07 V_low
+ 3.932010000e-07 V_low
+ 3.933000000e-07 V_low
+ 3.933010000e-07 V_low
+ 3.934000000e-07 V_low
+ 3.934010000e-07 V_low
+ 3.935000000e-07 V_low
+ 3.935010000e-07 V_low
+ 3.936000000e-07 V_low
+ 3.936010000e-07 V_low
+ 3.937000000e-07 V_low
+ 3.937010000e-07 V_low
+ 3.938000000e-07 V_low
+ 3.938010000e-07 V_low
+ 3.939000000e-07 V_low
+ 3.939010000e-07 V_low
+ 3.940000000e-07 V_low
+ 3.940010000e-07 V_low
+ 3.941000000e-07 V_low
+ 3.941010000e-07 V_low
+ 3.942000000e-07 V_low
+ 3.942010000e-07 V_low
+ 3.943000000e-07 V_low
+ 3.943010000e-07 V_low
+ 3.944000000e-07 V_low
+ 3.944010000e-07 V_low
+ 3.945000000e-07 V_low
+ 3.945010000e-07 V_low
+ 3.946000000e-07 V_low
+ 3.946010000e-07 V_low
+ 3.947000000e-07 V_low
+ 3.947010000e-07 V_low
+ 3.948000000e-07 V_low
+ 3.948010000e-07 V_low
+ 3.949000000e-07 V_low
+ 3.949010000e-07 V_low
+ 3.950000000e-07 V_low
+ 3.950010000e-07 V_low
+ 3.951000000e-07 V_low
+ 3.951010000e-07 V_low
+ 3.952000000e-07 V_low
+ 3.952010000e-07 V_low
+ 3.953000000e-07 V_low
+ 3.953010000e-07 V_low
+ 3.954000000e-07 V_low
+ 3.954010000e-07 V_low
+ 3.955000000e-07 V_low
+ 3.955010000e-07 V_low
+ 3.956000000e-07 V_low
+ 3.956010000e-07 V_low
+ 3.957000000e-07 V_low
+ 3.957010000e-07 V_low
+ 3.958000000e-07 V_low
+ 3.958010000e-07 V_low
+ 3.959000000e-07 V_low
+ 3.959010000e-07 V_low
+ 3.960000000e-07 V_low
+ 3.960010000e-07 V_low
+ 3.961000000e-07 V_low
+ 3.961010000e-07 V_low
+ 3.962000000e-07 V_low
+ 3.962010000e-07 V_low
+ 3.963000000e-07 V_low
+ 3.963010000e-07 V_low
+ 3.964000000e-07 V_low
+ 3.964010000e-07 V_low
+ 3.965000000e-07 V_low
+ 3.965010000e-07 V_low
+ 3.966000000e-07 V_low
+ 3.966010000e-07 V_low
+ 3.967000000e-07 V_low
+ 3.967010000e-07 V_low
+ 3.968000000e-07 V_low
+ 3.968010000e-07 V_low
+ 3.969000000e-07 V_low
+ 3.969010000e-07 V_low
+ 3.970000000e-07 V_low
+ 3.970010000e-07 V_low
+ 3.971000000e-07 V_low
+ 3.971010000e-07 V_low
+ 3.972000000e-07 V_low
+ 3.972010000e-07 V_low
+ 3.973000000e-07 V_low
+ 3.973010000e-07 V_low
+ 3.974000000e-07 V_low
+ 3.974010000e-07 V_low
+ 3.975000000e-07 V_low
+ 3.975010000e-07 V_low
+ 3.976000000e-07 V_low
+ 3.976010000e-07 V_low
+ 3.977000000e-07 V_low
+ 3.977010000e-07 V_low
+ 3.978000000e-07 V_low
+ 3.978010000e-07 V_low
+ 3.979000000e-07 V_low
+ 3.979010000e-07 V_low
+ 3.980000000e-07 V_low
+ 3.980010000e-07 V_low
+ 3.981000000e-07 V_low
+ 3.981010000e-07 V_low
+ 3.982000000e-07 V_low
+ 3.982010000e-07 V_low
+ 3.983000000e-07 V_low
+ 3.983010000e-07 V_low
+ 3.984000000e-07 V_low
+ 3.984010000e-07 V_low
+ 3.985000000e-07 V_low
+ 3.985010000e-07 V_low
+ 3.986000000e-07 V_low
+ 3.986010000e-07 V_low
+ 3.987000000e-07 V_low
+ 3.987010000e-07 V_low
+ 3.988000000e-07 V_low
+ 3.988010000e-07 V_low
+ 3.989000000e-07 V_low
+ 3.989010000e-07 V_low
+ 3.990000000e-07 V_low
+ 3.990010000e-07 V_low
+ 3.991000000e-07 V_low
+ 3.991010000e-07 V_low
+ 3.992000000e-07 V_low
+ 3.992010000e-07 V_low
+ 3.993000000e-07 V_low
+ 3.993010000e-07 V_low
+ 3.994000000e-07 V_low
+ 3.994010000e-07 V_low
+ 3.995000000e-07 V_low
+ 3.995010000e-07 V_low
+ 3.996000000e-07 V_low
+ 3.996010000e-07 V_low
+ 3.997000000e-07 V_low
+ 3.997010000e-07 V_low
+ 3.998000000e-07 V_low
+ 3.998010000e-07 V_low
+ 3.999000000e-07 V_low
+ 3.999010000e-07 V_hig
+ 4.000000000e-07 V_hig
+ 4.000010000e-07 V_hig
+ 4.001000000e-07 V_hig
+ 4.001010000e-07 V_hig
+ 4.002000000e-07 V_hig
+ 4.002010000e-07 V_hig
+ 4.003000000e-07 V_hig
+ 4.003010000e-07 V_hig
+ 4.004000000e-07 V_hig
+ 4.004010000e-07 V_hig
+ 4.005000000e-07 V_hig
+ 4.005010000e-07 V_hig
+ 4.006000000e-07 V_hig
+ 4.006010000e-07 V_hig
+ 4.007000000e-07 V_hig
+ 4.007010000e-07 V_hig
+ 4.008000000e-07 V_hig
+ 4.008010000e-07 V_hig
+ 4.009000000e-07 V_hig
+ 4.009010000e-07 V_low
+ 4.010000000e-07 V_low
+ 4.010010000e-07 V_low
+ 4.011000000e-07 V_low
+ 4.011010000e-07 V_low
+ 4.012000000e-07 V_low
+ 4.012010000e-07 V_low
+ 4.013000000e-07 V_low
+ 4.013010000e-07 V_low
+ 4.014000000e-07 V_low
+ 4.014010000e-07 V_low
+ 4.015000000e-07 V_low
+ 4.015010000e-07 V_low
+ 4.016000000e-07 V_low
+ 4.016010000e-07 V_low
+ 4.017000000e-07 V_low
+ 4.017010000e-07 V_low
+ 4.018000000e-07 V_low
+ 4.018010000e-07 V_low
+ 4.019000000e-07 V_low
+ 4.019010000e-07 V_hig
+ 4.020000000e-07 V_hig
+ 4.020010000e-07 V_hig
+ 4.021000000e-07 V_hig
+ 4.021010000e-07 V_hig
+ 4.022000000e-07 V_hig
+ 4.022010000e-07 V_hig
+ 4.023000000e-07 V_hig
+ 4.023010000e-07 V_hig
+ 4.024000000e-07 V_hig
+ 4.024010000e-07 V_hig
+ 4.025000000e-07 V_hig
+ 4.025010000e-07 V_hig
+ 4.026000000e-07 V_hig
+ 4.026010000e-07 V_hig
+ 4.027000000e-07 V_hig
+ 4.027010000e-07 V_hig
+ 4.028000000e-07 V_hig
+ 4.028010000e-07 V_hig
+ 4.029000000e-07 V_hig
+ 4.029010000e-07 V_low
+ 4.030000000e-07 V_low
+ 4.030010000e-07 V_low
+ 4.031000000e-07 V_low
+ 4.031010000e-07 V_low
+ 4.032000000e-07 V_low
+ 4.032010000e-07 V_low
+ 4.033000000e-07 V_low
+ 4.033010000e-07 V_low
+ 4.034000000e-07 V_low
+ 4.034010000e-07 V_low
+ 4.035000000e-07 V_low
+ 4.035010000e-07 V_low
+ 4.036000000e-07 V_low
+ 4.036010000e-07 V_low
+ 4.037000000e-07 V_low
+ 4.037010000e-07 V_low
+ 4.038000000e-07 V_low
+ 4.038010000e-07 V_low
+ 4.039000000e-07 V_low
+ 4.039010000e-07 V_hig
+ 4.040000000e-07 V_hig
+ 4.040010000e-07 V_hig
+ 4.041000000e-07 V_hig
+ 4.041010000e-07 V_hig
+ 4.042000000e-07 V_hig
+ 4.042010000e-07 V_hig
+ 4.043000000e-07 V_hig
+ 4.043010000e-07 V_hig
+ 4.044000000e-07 V_hig
+ 4.044010000e-07 V_hig
+ 4.045000000e-07 V_hig
+ 4.045010000e-07 V_hig
+ 4.046000000e-07 V_hig
+ 4.046010000e-07 V_hig
+ 4.047000000e-07 V_hig
+ 4.047010000e-07 V_hig
+ 4.048000000e-07 V_hig
+ 4.048010000e-07 V_hig
+ 4.049000000e-07 V_hig
+ 4.049010000e-07 V_low
+ 4.050000000e-07 V_low
+ 4.050010000e-07 V_low
+ 4.051000000e-07 V_low
+ 4.051010000e-07 V_low
+ 4.052000000e-07 V_low
+ 4.052010000e-07 V_low
+ 4.053000000e-07 V_low
+ 4.053010000e-07 V_low
+ 4.054000000e-07 V_low
+ 4.054010000e-07 V_low
+ 4.055000000e-07 V_low
+ 4.055010000e-07 V_low
+ 4.056000000e-07 V_low
+ 4.056010000e-07 V_low
+ 4.057000000e-07 V_low
+ 4.057010000e-07 V_low
+ 4.058000000e-07 V_low
+ 4.058010000e-07 V_low
+ 4.059000000e-07 V_low
+ 4.059010000e-07 V_low
+ 4.060000000e-07 V_low
+ 4.060010000e-07 V_low
+ 4.061000000e-07 V_low
+ 4.061010000e-07 V_low
+ 4.062000000e-07 V_low
+ 4.062010000e-07 V_low
+ 4.063000000e-07 V_low
+ 4.063010000e-07 V_low
+ 4.064000000e-07 V_low
+ 4.064010000e-07 V_low
+ 4.065000000e-07 V_low
+ 4.065010000e-07 V_low
+ 4.066000000e-07 V_low
+ 4.066010000e-07 V_low
+ 4.067000000e-07 V_low
+ 4.067010000e-07 V_low
+ 4.068000000e-07 V_low
+ 4.068010000e-07 V_low
+ 4.069000000e-07 V_low
+ 4.069010000e-07 V_low
+ 4.070000000e-07 V_low
+ 4.070010000e-07 V_low
+ 4.071000000e-07 V_low
+ 4.071010000e-07 V_low
+ 4.072000000e-07 V_low
+ 4.072010000e-07 V_low
+ 4.073000000e-07 V_low
+ 4.073010000e-07 V_low
+ 4.074000000e-07 V_low
+ 4.074010000e-07 V_low
+ 4.075000000e-07 V_low
+ 4.075010000e-07 V_low
+ 4.076000000e-07 V_low
+ 4.076010000e-07 V_low
+ 4.077000000e-07 V_low
+ 4.077010000e-07 V_low
+ 4.078000000e-07 V_low
+ 4.078010000e-07 V_low
+ 4.079000000e-07 V_low
+ 4.079010000e-07 V_low
+ 4.080000000e-07 V_low
+ 4.080010000e-07 V_low
+ 4.081000000e-07 V_low
+ 4.081010000e-07 V_low
+ 4.082000000e-07 V_low
+ 4.082010000e-07 V_low
+ 4.083000000e-07 V_low
+ 4.083010000e-07 V_low
+ 4.084000000e-07 V_low
+ 4.084010000e-07 V_low
+ 4.085000000e-07 V_low
+ 4.085010000e-07 V_low
+ 4.086000000e-07 V_low
+ 4.086010000e-07 V_low
+ 4.087000000e-07 V_low
+ 4.087010000e-07 V_low
+ 4.088000000e-07 V_low
+ 4.088010000e-07 V_low
+ 4.089000000e-07 V_low
+ 4.089010000e-07 V_hig
+ 4.090000000e-07 V_hig
+ 4.090010000e-07 V_hig
+ 4.091000000e-07 V_hig
+ 4.091010000e-07 V_hig
+ 4.092000000e-07 V_hig
+ 4.092010000e-07 V_hig
+ 4.093000000e-07 V_hig
+ 4.093010000e-07 V_hig
+ 4.094000000e-07 V_hig
+ 4.094010000e-07 V_hig
+ 4.095000000e-07 V_hig
+ 4.095010000e-07 V_hig
+ 4.096000000e-07 V_hig
+ 4.096010000e-07 V_hig
+ 4.097000000e-07 V_hig
+ 4.097010000e-07 V_hig
+ 4.098000000e-07 V_hig
+ 4.098010000e-07 V_hig
+ 4.099000000e-07 V_hig
+ 4.099010000e-07 V_hig
+ 4.100000000e-07 V_hig
+ 4.100010000e-07 V_hig
+ 4.101000000e-07 V_hig
+ 4.101010000e-07 V_hig
+ 4.102000000e-07 V_hig
+ 4.102010000e-07 V_hig
+ 4.103000000e-07 V_hig
+ 4.103010000e-07 V_hig
+ 4.104000000e-07 V_hig
+ 4.104010000e-07 V_hig
+ 4.105000000e-07 V_hig
+ 4.105010000e-07 V_hig
+ 4.106000000e-07 V_hig
+ 4.106010000e-07 V_hig
+ 4.107000000e-07 V_hig
+ 4.107010000e-07 V_hig
+ 4.108000000e-07 V_hig
+ 4.108010000e-07 V_hig
+ 4.109000000e-07 V_hig
+ 4.109010000e-07 V_low
+ 4.110000000e-07 V_low
+ 4.110010000e-07 V_low
+ 4.111000000e-07 V_low
+ 4.111010000e-07 V_low
+ 4.112000000e-07 V_low
+ 4.112010000e-07 V_low
+ 4.113000000e-07 V_low
+ 4.113010000e-07 V_low
+ 4.114000000e-07 V_low
+ 4.114010000e-07 V_low
+ 4.115000000e-07 V_low
+ 4.115010000e-07 V_low
+ 4.116000000e-07 V_low
+ 4.116010000e-07 V_low
+ 4.117000000e-07 V_low
+ 4.117010000e-07 V_low
+ 4.118000000e-07 V_low
+ 4.118010000e-07 V_low
+ 4.119000000e-07 V_low
+ 4.119010000e-07 V_low
+ 4.120000000e-07 V_low
+ 4.120010000e-07 V_low
+ 4.121000000e-07 V_low
+ 4.121010000e-07 V_low
+ 4.122000000e-07 V_low
+ 4.122010000e-07 V_low
+ 4.123000000e-07 V_low
+ 4.123010000e-07 V_low
+ 4.124000000e-07 V_low
+ 4.124010000e-07 V_low
+ 4.125000000e-07 V_low
+ 4.125010000e-07 V_low
+ 4.126000000e-07 V_low
+ 4.126010000e-07 V_low
+ 4.127000000e-07 V_low
+ 4.127010000e-07 V_low
+ 4.128000000e-07 V_low
+ 4.128010000e-07 V_low
+ 4.129000000e-07 V_low
+ 4.129010000e-07 V_hig
+ 4.130000000e-07 V_hig
+ 4.130010000e-07 V_hig
+ 4.131000000e-07 V_hig
+ 4.131010000e-07 V_hig
+ 4.132000000e-07 V_hig
+ 4.132010000e-07 V_hig
+ 4.133000000e-07 V_hig
+ 4.133010000e-07 V_hig
+ 4.134000000e-07 V_hig
+ 4.134010000e-07 V_hig
+ 4.135000000e-07 V_hig
+ 4.135010000e-07 V_hig
+ 4.136000000e-07 V_hig
+ 4.136010000e-07 V_hig
+ 4.137000000e-07 V_hig
+ 4.137010000e-07 V_hig
+ 4.138000000e-07 V_hig
+ 4.138010000e-07 V_hig
+ 4.139000000e-07 V_hig
+ 4.139010000e-07 V_hig
+ 4.140000000e-07 V_hig
+ 4.140010000e-07 V_hig
+ 4.141000000e-07 V_hig
+ 4.141010000e-07 V_hig
+ 4.142000000e-07 V_hig
+ 4.142010000e-07 V_hig
+ 4.143000000e-07 V_hig
+ 4.143010000e-07 V_hig
+ 4.144000000e-07 V_hig
+ 4.144010000e-07 V_hig
+ 4.145000000e-07 V_hig
+ 4.145010000e-07 V_hig
+ 4.146000000e-07 V_hig
+ 4.146010000e-07 V_hig
+ 4.147000000e-07 V_hig
+ 4.147010000e-07 V_hig
+ 4.148000000e-07 V_hig
+ 4.148010000e-07 V_hig
+ 4.149000000e-07 V_hig
+ 4.149010000e-07 V_low
+ 4.150000000e-07 V_low
+ 4.150010000e-07 V_low
+ 4.151000000e-07 V_low
+ 4.151010000e-07 V_low
+ 4.152000000e-07 V_low
+ 4.152010000e-07 V_low
+ 4.153000000e-07 V_low
+ 4.153010000e-07 V_low
+ 4.154000000e-07 V_low
+ 4.154010000e-07 V_low
+ 4.155000000e-07 V_low
+ 4.155010000e-07 V_low
+ 4.156000000e-07 V_low
+ 4.156010000e-07 V_low
+ 4.157000000e-07 V_low
+ 4.157010000e-07 V_low
+ 4.158000000e-07 V_low
+ 4.158010000e-07 V_low
+ 4.159000000e-07 V_low
+ 4.159010000e-07 V_low
+ 4.160000000e-07 V_low
+ 4.160010000e-07 V_low
+ 4.161000000e-07 V_low
+ 4.161010000e-07 V_low
+ 4.162000000e-07 V_low
+ 4.162010000e-07 V_low
+ 4.163000000e-07 V_low
+ 4.163010000e-07 V_low
+ 4.164000000e-07 V_low
+ 4.164010000e-07 V_low
+ 4.165000000e-07 V_low
+ 4.165010000e-07 V_low
+ 4.166000000e-07 V_low
+ 4.166010000e-07 V_low
+ 4.167000000e-07 V_low
+ 4.167010000e-07 V_low
+ 4.168000000e-07 V_low
+ 4.168010000e-07 V_low
+ 4.169000000e-07 V_low
+ 4.169010000e-07 V_low
+ 4.170000000e-07 V_low
+ 4.170010000e-07 V_low
+ 4.171000000e-07 V_low
+ 4.171010000e-07 V_low
+ 4.172000000e-07 V_low
+ 4.172010000e-07 V_low
+ 4.173000000e-07 V_low
+ 4.173010000e-07 V_low
+ 4.174000000e-07 V_low
+ 4.174010000e-07 V_low
+ 4.175000000e-07 V_low
+ 4.175010000e-07 V_low
+ 4.176000000e-07 V_low
+ 4.176010000e-07 V_low
+ 4.177000000e-07 V_low
+ 4.177010000e-07 V_low
+ 4.178000000e-07 V_low
+ 4.178010000e-07 V_low
+ 4.179000000e-07 V_low
+ 4.179010000e-07 V_low
+ 4.180000000e-07 V_low
+ 4.180010000e-07 V_low
+ 4.181000000e-07 V_low
+ 4.181010000e-07 V_low
+ 4.182000000e-07 V_low
+ 4.182010000e-07 V_low
+ 4.183000000e-07 V_low
+ 4.183010000e-07 V_low
+ 4.184000000e-07 V_low
+ 4.184010000e-07 V_low
+ 4.185000000e-07 V_low
+ 4.185010000e-07 V_low
+ 4.186000000e-07 V_low
+ 4.186010000e-07 V_low
+ 4.187000000e-07 V_low
+ 4.187010000e-07 V_low
+ 4.188000000e-07 V_low
+ 4.188010000e-07 V_low
+ 4.189000000e-07 V_low
+ 4.189010000e-07 V_hig
+ 4.190000000e-07 V_hig
+ 4.190010000e-07 V_hig
+ 4.191000000e-07 V_hig
+ 4.191010000e-07 V_hig
+ 4.192000000e-07 V_hig
+ 4.192010000e-07 V_hig
+ 4.193000000e-07 V_hig
+ 4.193010000e-07 V_hig
+ 4.194000000e-07 V_hig
+ 4.194010000e-07 V_hig
+ 4.195000000e-07 V_hig
+ 4.195010000e-07 V_hig
+ 4.196000000e-07 V_hig
+ 4.196010000e-07 V_hig
+ 4.197000000e-07 V_hig
+ 4.197010000e-07 V_hig
+ 4.198000000e-07 V_hig
+ 4.198010000e-07 V_hig
+ 4.199000000e-07 V_hig
+ 4.199010000e-07 V_low
+ 4.200000000e-07 V_low
+ 4.200010000e-07 V_low
+ 4.201000000e-07 V_low
+ 4.201010000e-07 V_low
+ 4.202000000e-07 V_low
+ 4.202010000e-07 V_low
+ 4.203000000e-07 V_low
+ 4.203010000e-07 V_low
+ 4.204000000e-07 V_low
+ 4.204010000e-07 V_low
+ 4.205000000e-07 V_low
+ 4.205010000e-07 V_low
+ 4.206000000e-07 V_low
+ 4.206010000e-07 V_low
+ 4.207000000e-07 V_low
+ 4.207010000e-07 V_low
+ 4.208000000e-07 V_low
+ 4.208010000e-07 V_low
+ 4.209000000e-07 V_low
+ 4.209010000e-07 V_low
+ 4.210000000e-07 V_low
+ 4.210010000e-07 V_low
+ 4.211000000e-07 V_low
+ 4.211010000e-07 V_low
+ 4.212000000e-07 V_low
+ 4.212010000e-07 V_low
+ 4.213000000e-07 V_low
+ 4.213010000e-07 V_low
+ 4.214000000e-07 V_low
+ 4.214010000e-07 V_low
+ 4.215000000e-07 V_low
+ 4.215010000e-07 V_low
+ 4.216000000e-07 V_low
+ 4.216010000e-07 V_low
+ 4.217000000e-07 V_low
+ 4.217010000e-07 V_low
+ 4.218000000e-07 V_low
+ 4.218010000e-07 V_low
+ 4.219000000e-07 V_low
+ 4.219010000e-07 V_low
+ 4.220000000e-07 V_low
+ 4.220010000e-07 V_low
+ 4.221000000e-07 V_low
+ 4.221010000e-07 V_low
+ 4.222000000e-07 V_low
+ 4.222010000e-07 V_low
+ 4.223000000e-07 V_low
+ 4.223010000e-07 V_low
+ 4.224000000e-07 V_low
+ 4.224010000e-07 V_low
+ 4.225000000e-07 V_low
+ 4.225010000e-07 V_low
+ 4.226000000e-07 V_low
+ 4.226010000e-07 V_low
+ 4.227000000e-07 V_low
+ 4.227010000e-07 V_low
+ 4.228000000e-07 V_low
+ 4.228010000e-07 V_low
+ 4.229000000e-07 V_low
+ 4.229010000e-07 V_low
+ 4.230000000e-07 V_low
+ 4.230010000e-07 V_low
+ 4.231000000e-07 V_low
+ 4.231010000e-07 V_low
+ 4.232000000e-07 V_low
+ 4.232010000e-07 V_low
+ 4.233000000e-07 V_low
+ 4.233010000e-07 V_low
+ 4.234000000e-07 V_low
+ 4.234010000e-07 V_low
+ 4.235000000e-07 V_low
+ 4.235010000e-07 V_low
+ 4.236000000e-07 V_low
+ 4.236010000e-07 V_low
+ 4.237000000e-07 V_low
+ 4.237010000e-07 V_low
+ 4.238000000e-07 V_low
+ 4.238010000e-07 V_low
+ 4.239000000e-07 V_low
+ 4.239010000e-07 V_low
+ 4.240000000e-07 V_low
+ 4.240010000e-07 V_low
+ 4.241000000e-07 V_low
+ 4.241010000e-07 V_low
+ 4.242000000e-07 V_low
+ 4.242010000e-07 V_low
+ 4.243000000e-07 V_low
+ 4.243010000e-07 V_low
+ 4.244000000e-07 V_low
+ 4.244010000e-07 V_low
+ 4.245000000e-07 V_low
+ 4.245010000e-07 V_low
+ 4.246000000e-07 V_low
+ 4.246010000e-07 V_low
+ 4.247000000e-07 V_low
+ 4.247010000e-07 V_low
+ 4.248000000e-07 V_low
+ 4.248010000e-07 V_low
+ 4.249000000e-07 V_low
+ 4.249010000e-07 V_low
+ 4.250000000e-07 V_low
+ 4.250010000e-07 V_low
+ 4.251000000e-07 V_low
+ 4.251010000e-07 V_low
+ 4.252000000e-07 V_low
+ 4.252010000e-07 V_low
+ 4.253000000e-07 V_low
+ 4.253010000e-07 V_low
+ 4.254000000e-07 V_low
+ 4.254010000e-07 V_low
+ 4.255000000e-07 V_low
+ 4.255010000e-07 V_low
+ 4.256000000e-07 V_low
+ 4.256010000e-07 V_low
+ 4.257000000e-07 V_low
+ 4.257010000e-07 V_low
+ 4.258000000e-07 V_low
+ 4.258010000e-07 V_low
+ 4.259000000e-07 V_low
+ 4.259010000e-07 V_hig
+ 4.260000000e-07 V_hig
+ 4.260010000e-07 V_hig
+ 4.261000000e-07 V_hig
+ 4.261010000e-07 V_hig
+ 4.262000000e-07 V_hig
+ 4.262010000e-07 V_hig
+ 4.263000000e-07 V_hig
+ 4.263010000e-07 V_hig
+ 4.264000000e-07 V_hig
+ 4.264010000e-07 V_hig
+ 4.265000000e-07 V_hig
+ 4.265010000e-07 V_hig
+ 4.266000000e-07 V_hig
+ 4.266010000e-07 V_hig
+ 4.267000000e-07 V_hig
+ 4.267010000e-07 V_hig
+ 4.268000000e-07 V_hig
+ 4.268010000e-07 V_hig
+ 4.269000000e-07 V_hig
+ 4.269010000e-07 V_hig
+ 4.270000000e-07 V_hig
+ 4.270010000e-07 V_hig
+ 4.271000000e-07 V_hig
+ 4.271010000e-07 V_hig
+ 4.272000000e-07 V_hig
+ 4.272010000e-07 V_hig
+ 4.273000000e-07 V_hig
+ 4.273010000e-07 V_hig
+ 4.274000000e-07 V_hig
+ 4.274010000e-07 V_hig
+ 4.275000000e-07 V_hig
+ 4.275010000e-07 V_hig
+ 4.276000000e-07 V_hig
+ 4.276010000e-07 V_hig
+ 4.277000000e-07 V_hig
+ 4.277010000e-07 V_hig
+ 4.278000000e-07 V_hig
+ 4.278010000e-07 V_hig
+ 4.279000000e-07 V_hig
+ 4.279010000e-07 V_low
+ 4.280000000e-07 V_low
+ 4.280010000e-07 V_low
+ 4.281000000e-07 V_low
+ 4.281010000e-07 V_low
+ 4.282000000e-07 V_low
+ 4.282010000e-07 V_low
+ 4.283000000e-07 V_low
+ 4.283010000e-07 V_low
+ 4.284000000e-07 V_low
+ 4.284010000e-07 V_low
+ 4.285000000e-07 V_low
+ 4.285010000e-07 V_low
+ 4.286000000e-07 V_low
+ 4.286010000e-07 V_low
+ 4.287000000e-07 V_low
+ 4.287010000e-07 V_low
+ 4.288000000e-07 V_low
+ 4.288010000e-07 V_low
+ 4.289000000e-07 V_low
+ 4.289010000e-07 V_hig
+ 4.290000000e-07 V_hig
+ 4.290010000e-07 V_hig
+ 4.291000000e-07 V_hig
+ 4.291010000e-07 V_hig
+ 4.292000000e-07 V_hig
+ 4.292010000e-07 V_hig
+ 4.293000000e-07 V_hig
+ 4.293010000e-07 V_hig
+ 4.294000000e-07 V_hig
+ 4.294010000e-07 V_hig
+ 4.295000000e-07 V_hig
+ 4.295010000e-07 V_hig
+ 4.296000000e-07 V_hig
+ 4.296010000e-07 V_hig
+ 4.297000000e-07 V_hig
+ 4.297010000e-07 V_hig
+ 4.298000000e-07 V_hig
+ 4.298010000e-07 V_hig
+ 4.299000000e-07 V_hig
+ 4.299010000e-07 V_hig
+ 4.300000000e-07 V_hig
+ 4.300010000e-07 V_hig
+ 4.301000000e-07 V_hig
+ 4.301010000e-07 V_hig
+ 4.302000000e-07 V_hig
+ 4.302010000e-07 V_hig
+ 4.303000000e-07 V_hig
+ 4.303010000e-07 V_hig
+ 4.304000000e-07 V_hig
+ 4.304010000e-07 V_hig
+ 4.305000000e-07 V_hig
+ 4.305010000e-07 V_hig
+ 4.306000000e-07 V_hig
+ 4.306010000e-07 V_hig
+ 4.307000000e-07 V_hig
+ 4.307010000e-07 V_hig
+ 4.308000000e-07 V_hig
+ 4.308010000e-07 V_hig
+ 4.309000000e-07 V_hig
+ 4.309010000e-07 V_low
+ 4.310000000e-07 V_low
+ 4.310010000e-07 V_low
+ 4.311000000e-07 V_low
+ 4.311010000e-07 V_low
+ 4.312000000e-07 V_low
+ 4.312010000e-07 V_low
+ 4.313000000e-07 V_low
+ 4.313010000e-07 V_low
+ 4.314000000e-07 V_low
+ 4.314010000e-07 V_low
+ 4.315000000e-07 V_low
+ 4.315010000e-07 V_low
+ 4.316000000e-07 V_low
+ 4.316010000e-07 V_low
+ 4.317000000e-07 V_low
+ 4.317010000e-07 V_low
+ 4.318000000e-07 V_low
+ 4.318010000e-07 V_low
+ 4.319000000e-07 V_low
+ 4.319010000e-07 V_hig
+ 4.320000000e-07 V_hig
+ 4.320010000e-07 V_hig
+ 4.321000000e-07 V_hig
+ 4.321010000e-07 V_hig
+ 4.322000000e-07 V_hig
+ 4.322010000e-07 V_hig
+ 4.323000000e-07 V_hig
+ 4.323010000e-07 V_hig
+ 4.324000000e-07 V_hig
+ 4.324010000e-07 V_hig
+ 4.325000000e-07 V_hig
+ 4.325010000e-07 V_hig
+ 4.326000000e-07 V_hig
+ 4.326010000e-07 V_hig
+ 4.327000000e-07 V_hig
+ 4.327010000e-07 V_hig
+ 4.328000000e-07 V_hig
+ 4.328010000e-07 V_hig
+ 4.329000000e-07 V_hig
+ 4.329010000e-07 V_hig
+ 4.330000000e-07 V_hig
+ 4.330010000e-07 V_hig
+ 4.331000000e-07 V_hig
+ 4.331010000e-07 V_hig
+ 4.332000000e-07 V_hig
+ 4.332010000e-07 V_hig
+ 4.333000000e-07 V_hig
+ 4.333010000e-07 V_hig
+ 4.334000000e-07 V_hig
+ 4.334010000e-07 V_hig
+ 4.335000000e-07 V_hig
+ 4.335010000e-07 V_hig
+ 4.336000000e-07 V_hig
+ 4.336010000e-07 V_hig
+ 4.337000000e-07 V_hig
+ 4.337010000e-07 V_hig
+ 4.338000000e-07 V_hig
+ 4.338010000e-07 V_hig
+ 4.339000000e-07 V_hig
+ 4.339010000e-07 V_hig
+ 4.340000000e-07 V_hig
+ 4.340010000e-07 V_hig
+ 4.341000000e-07 V_hig
+ 4.341010000e-07 V_hig
+ 4.342000000e-07 V_hig
+ 4.342010000e-07 V_hig
+ 4.343000000e-07 V_hig
+ 4.343010000e-07 V_hig
+ 4.344000000e-07 V_hig
+ 4.344010000e-07 V_hig
+ 4.345000000e-07 V_hig
+ 4.345010000e-07 V_hig
+ 4.346000000e-07 V_hig
+ 4.346010000e-07 V_hig
+ 4.347000000e-07 V_hig
+ 4.347010000e-07 V_hig
+ 4.348000000e-07 V_hig
+ 4.348010000e-07 V_hig
+ 4.349000000e-07 V_hig
+ 4.349010000e-07 V_hig
+ 4.350000000e-07 V_hig
+ 4.350010000e-07 V_hig
+ 4.351000000e-07 V_hig
+ 4.351010000e-07 V_hig
+ 4.352000000e-07 V_hig
+ 4.352010000e-07 V_hig
+ 4.353000000e-07 V_hig
+ 4.353010000e-07 V_hig
+ 4.354000000e-07 V_hig
+ 4.354010000e-07 V_hig
+ 4.355000000e-07 V_hig
+ 4.355010000e-07 V_hig
+ 4.356000000e-07 V_hig
+ 4.356010000e-07 V_hig
+ 4.357000000e-07 V_hig
+ 4.357010000e-07 V_hig
+ 4.358000000e-07 V_hig
+ 4.358010000e-07 V_hig
+ 4.359000000e-07 V_hig
+ 4.359010000e-07 V_low
+ 4.360000000e-07 V_low
+ 4.360010000e-07 V_low
+ 4.361000000e-07 V_low
+ 4.361010000e-07 V_low
+ 4.362000000e-07 V_low
+ 4.362010000e-07 V_low
+ 4.363000000e-07 V_low
+ 4.363010000e-07 V_low
+ 4.364000000e-07 V_low
+ 4.364010000e-07 V_low
+ 4.365000000e-07 V_low
+ 4.365010000e-07 V_low
+ 4.366000000e-07 V_low
+ 4.366010000e-07 V_low
+ 4.367000000e-07 V_low
+ 4.367010000e-07 V_low
+ 4.368000000e-07 V_low
+ 4.368010000e-07 V_low
+ 4.369000000e-07 V_low
+ 4.369010000e-07 V_hig
+ 4.370000000e-07 V_hig
+ 4.370010000e-07 V_hig
+ 4.371000000e-07 V_hig
+ 4.371010000e-07 V_hig
+ 4.372000000e-07 V_hig
+ 4.372010000e-07 V_hig
+ 4.373000000e-07 V_hig
+ 4.373010000e-07 V_hig
+ 4.374000000e-07 V_hig
+ 4.374010000e-07 V_hig
+ 4.375000000e-07 V_hig
+ 4.375010000e-07 V_hig
+ 4.376000000e-07 V_hig
+ 4.376010000e-07 V_hig
+ 4.377000000e-07 V_hig
+ 4.377010000e-07 V_hig
+ 4.378000000e-07 V_hig
+ 4.378010000e-07 V_hig
+ 4.379000000e-07 V_hig
+ 4.379010000e-07 V_hig
+ 4.380000000e-07 V_hig
+ 4.380010000e-07 V_hig
+ 4.381000000e-07 V_hig
+ 4.381010000e-07 V_hig
+ 4.382000000e-07 V_hig
+ 4.382010000e-07 V_hig
+ 4.383000000e-07 V_hig
+ 4.383010000e-07 V_hig
+ 4.384000000e-07 V_hig
+ 4.384010000e-07 V_hig
+ 4.385000000e-07 V_hig
+ 4.385010000e-07 V_hig
+ 4.386000000e-07 V_hig
+ 4.386010000e-07 V_hig
+ 4.387000000e-07 V_hig
+ 4.387010000e-07 V_hig
+ 4.388000000e-07 V_hig
+ 4.388010000e-07 V_hig
+ 4.389000000e-07 V_hig
+ 4.389010000e-07 V_hig
+ 4.390000000e-07 V_hig
+ 4.390010000e-07 V_hig
+ 4.391000000e-07 V_hig
+ 4.391010000e-07 V_hig
+ 4.392000000e-07 V_hig
+ 4.392010000e-07 V_hig
+ 4.393000000e-07 V_hig
+ 4.393010000e-07 V_hig
+ 4.394000000e-07 V_hig
+ 4.394010000e-07 V_hig
+ 4.395000000e-07 V_hig
+ 4.395010000e-07 V_hig
+ 4.396000000e-07 V_hig
+ 4.396010000e-07 V_hig
+ 4.397000000e-07 V_hig
+ 4.397010000e-07 V_hig
+ 4.398000000e-07 V_hig
+ 4.398010000e-07 V_hig
+ 4.399000000e-07 V_hig
+ 4.399010000e-07 V_hig
+ 4.400000000e-07 V_hig
+ 4.400010000e-07 V_hig
+ 4.401000000e-07 V_hig
+ 4.401010000e-07 V_hig
+ 4.402000000e-07 V_hig
+ 4.402010000e-07 V_hig
+ 4.403000000e-07 V_hig
+ 4.403010000e-07 V_hig
+ 4.404000000e-07 V_hig
+ 4.404010000e-07 V_hig
+ 4.405000000e-07 V_hig
+ 4.405010000e-07 V_hig
+ 4.406000000e-07 V_hig
+ 4.406010000e-07 V_hig
+ 4.407000000e-07 V_hig
+ 4.407010000e-07 V_hig
+ 4.408000000e-07 V_hig
+ 4.408010000e-07 V_hig
+ 4.409000000e-07 V_hig
+ 4.409010000e-07 V_low
+ 4.410000000e-07 V_low
+ 4.410010000e-07 V_low
+ 4.411000000e-07 V_low
+ 4.411010000e-07 V_low
+ 4.412000000e-07 V_low
+ 4.412010000e-07 V_low
+ 4.413000000e-07 V_low
+ 4.413010000e-07 V_low
+ 4.414000000e-07 V_low
+ 4.414010000e-07 V_low
+ 4.415000000e-07 V_low
+ 4.415010000e-07 V_low
+ 4.416000000e-07 V_low
+ 4.416010000e-07 V_low
+ 4.417000000e-07 V_low
+ 4.417010000e-07 V_low
+ 4.418000000e-07 V_low
+ 4.418010000e-07 V_low
+ 4.419000000e-07 V_low
+ 4.419010000e-07 V_low
+ 4.420000000e-07 V_low
+ 4.420010000e-07 V_low
+ 4.421000000e-07 V_low
+ 4.421010000e-07 V_low
+ 4.422000000e-07 V_low
+ 4.422010000e-07 V_low
+ 4.423000000e-07 V_low
+ 4.423010000e-07 V_low
+ 4.424000000e-07 V_low
+ 4.424010000e-07 V_low
+ 4.425000000e-07 V_low
+ 4.425010000e-07 V_low
+ 4.426000000e-07 V_low
+ 4.426010000e-07 V_low
+ 4.427000000e-07 V_low
+ 4.427010000e-07 V_low
+ 4.428000000e-07 V_low
+ 4.428010000e-07 V_low
+ 4.429000000e-07 V_low
+ 4.429010000e-07 V_low
+ 4.430000000e-07 V_low
+ 4.430010000e-07 V_low
+ 4.431000000e-07 V_low
+ 4.431010000e-07 V_low
+ 4.432000000e-07 V_low
+ 4.432010000e-07 V_low
+ 4.433000000e-07 V_low
+ 4.433010000e-07 V_low
+ 4.434000000e-07 V_low
+ 4.434010000e-07 V_low
+ 4.435000000e-07 V_low
+ 4.435010000e-07 V_low
+ 4.436000000e-07 V_low
+ 4.436010000e-07 V_low
+ 4.437000000e-07 V_low
+ 4.437010000e-07 V_low
+ 4.438000000e-07 V_low
+ 4.438010000e-07 V_low
+ 4.439000000e-07 V_low
+ 4.439010000e-07 V_low
+ 4.440000000e-07 V_low
+ 4.440010000e-07 V_low
+ 4.441000000e-07 V_low
+ 4.441010000e-07 V_low
+ 4.442000000e-07 V_low
+ 4.442010000e-07 V_low
+ 4.443000000e-07 V_low
+ 4.443010000e-07 V_low
+ 4.444000000e-07 V_low
+ 4.444010000e-07 V_low
+ 4.445000000e-07 V_low
+ 4.445010000e-07 V_low
+ 4.446000000e-07 V_low
+ 4.446010000e-07 V_low
+ 4.447000000e-07 V_low
+ 4.447010000e-07 V_low
+ 4.448000000e-07 V_low
+ 4.448010000e-07 V_low
+ 4.449000000e-07 V_low
+ 4.449010000e-07 V_low
+ 4.450000000e-07 V_low
+ 4.450010000e-07 V_low
+ 4.451000000e-07 V_low
+ 4.451010000e-07 V_low
+ 4.452000000e-07 V_low
+ 4.452010000e-07 V_low
+ 4.453000000e-07 V_low
+ 4.453010000e-07 V_low
+ 4.454000000e-07 V_low
+ 4.454010000e-07 V_low
+ 4.455000000e-07 V_low
+ 4.455010000e-07 V_low
+ 4.456000000e-07 V_low
+ 4.456010000e-07 V_low
+ 4.457000000e-07 V_low
+ 4.457010000e-07 V_low
+ 4.458000000e-07 V_low
+ 4.458010000e-07 V_low
+ 4.459000000e-07 V_low
+ 4.459010000e-07 V_hig
+ 4.460000000e-07 V_hig
+ 4.460010000e-07 V_hig
+ 4.461000000e-07 V_hig
+ 4.461010000e-07 V_hig
+ 4.462000000e-07 V_hig
+ 4.462010000e-07 V_hig
+ 4.463000000e-07 V_hig
+ 4.463010000e-07 V_hig
+ 4.464000000e-07 V_hig
+ 4.464010000e-07 V_hig
+ 4.465000000e-07 V_hig
+ 4.465010000e-07 V_hig
+ 4.466000000e-07 V_hig
+ 4.466010000e-07 V_hig
+ 4.467000000e-07 V_hig
+ 4.467010000e-07 V_hig
+ 4.468000000e-07 V_hig
+ 4.468010000e-07 V_hig
+ 4.469000000e-07 V_hig
+ 4.469010000e-07 V_low
+ 4.470000000e-07 V_low
+ 4.470010000e-07 V_low
+ 4.471000000e-07 V_low
+ 4.471010000e-07 V_low
+ 4.472000000e-07 V_low
+ 4.472010000e-07 V_low
+ 4.473000000e-07 V_low
+ 4.473010000e-07 V_low
+ 4.474000000e-07 V_low
+ 4.474010000e-07 V_low
+ 4.475000000e-07 V_low
+ 4.475010000e-07 V_low
+ 4.476000000e-07 V_low
+ 4.476010000e-07 V_low
+ 4.477000000e-07 V_low
+ 4.477010000e-07 V_low
+ 4.478000000e-07 V_low
+ 4.478010000e-07 V_low
+ 4.479000000e-07 V_low
+ 4.479010000e-07 V_hig
+ 4.480000000e-07 V_hig
+ 4.480010000e-07 V_hig
+ 4.481000000e-07 V_hig
+ 4.481010000e-07 V_hig
+ 4.482000000e-07 V_hig
+ 4.482010000e-07 V_hig
+ 4.483000000e-07 V_hig
+ 4.483010000e-07 V_hig
+ 4.484000000e-07 V_hig
+ 4.484010000e-07 V_hig
+ 4.485000000e-07 V_hig
+ 4.485010000e-07 V_hig
+ 4.486000000e-07 V_hig
+ 4.486010000e-07 V_hig
+ 4.487000000e-07 V_hig
+ 4.487010000e-07 V_hig
+ 4.488000000e-07 V_hig
+ 4.488010000e-07 V_hig
+ 4.489000000e-07 V_hig
+ 4.489010000e-07 V_low
+ 4.490000000e-07 V_low
+ 4.490010000e-07 V_low
+ 4.491000000e-07 V_low
+ 4.491010000e-07 V_low
+ 4.492000000e-07 V_low
+ 4.492010000e-07 V_low
+ 4.493000000e-07 V_low
+ 4.493010000e-07 V_low
+ 4.494000000e-07 V_low
+ 4.494010000e-07 V_low
+ 4.495000000e-07 V_low
+ 4.495010000e-07 V_low
+ 4.496000000e-07 V_low
+ 4.496010000e-07 V_low
+ 4.497000000e-07 V_low
+ 4.497010000e-07 V_low
+ 4.498000000e-07 V_low
+ 4.498010000e-07 V_low
+ 4.499000000e-07 V_low
+ 4.499010000e-07 V_hig
+ 4.500000000e-07 V_hig
+ 4.500010000e-07 V_hig
+ 4.501000000e-07 V_hig
+ 4.501010000e-07 V_hig
+ 4.502000000e-07 V_hig
+ 4.502010000e-07 V_hig
+ 4.503000000e-07 V_hig
+ 4.503010000e-07 V_hig
+ 4.504000000e-07 V_hig
+ 4.504010000e-07 V_hig
+ 4.505000000e-07 V_hig
+ 4.505010000e-07 V_hig
+ 4.506000000e-07 V_hig
+ 4.506010000e-07 V_hig
+ 4.507000000e-07 V_hig
+ 4.507010000e-07 V_hig
+ 4.508000000e-07 V_hig
+ 4.508010000e-07 V_hig
+ 4.509000000e-07 V_hig
+ 4.509010000e-07 V_hig
+ 4.510000000e-07 V_hig
+ 4.510010000e-07 V_hig
+ 4.511000000e-07 V_hig
+ 4.511010000e-07 V_hig
+ 4.512000000e-07 V_hig
+ 4.512010000e-07 V_hig
+ 4.513000000e-07 V_hig
+ 4.513010000e-07 V_hig
+ 4.514000000e-07 V_hig
+ 4.514010000e-07 V_hig
+ 4.515000000e-07 V_hig
+ 4.515010000e-07 V_hig
+ 4.516000000e-07 V_hig
+ 4.516010000e-07 V_hig
+ 4.517000000e-07 V_hig
+ 4.517010000e-07 V_hig
+ 4.518000000e-07 V_hig
+ 4.518010000e-07 V_hig
+ 4.519000000e-07 V_hig
+ 4.519010000e-07 V_hig
+ 4.520000000e-07 V_hig
+ 4.520010000e-07 V_hig
+ 4.521000000e-07 V_hig
+ 4.521010000e-07 V_hig
+ 4.522000000e-07 V_hig
+ 4.522010000e-07 V_hig
+ 4.523000000e-07 V_hig
+ 4.523010000e-07 V_hig
+ 4.524000000e-07 V_hig
+ 4.524010000e-07 V_hig
+ 4.525000000e-07 V_hig
+ 4.525010000e-07 V_hig
+ 4.526000000e-07 V_hig
+ 4.526010000e-07 V_hig
+ 4.527000000e-07 V_hig
+ 4.527010000e-07 V_hig
+ 4.528000000e-07 V_hig
+ 4.528010000e-07 V_hig
+ 4.529000000e-07 V_hig
+ 4.529010000e-07 V_low
+ 4.530000000e-07 V_low
+ 4.530010000e-07 V_low
+ 4.531000000e-07 V_low
+ 4.531010000e-07 V_low
+ 4.532000000e-07 V_low
+ 4.532010000e-07 V_low
+ 4.533000000e-07 V_low
+ 4.533010000e-07 V_low
+ 4.534000000e-07 V_low
+ 4.534010000e-07 V_low
+ 4.535000000e-07 V_low
+ 4.535010000e-07 V_low
+ 4.536000000e-07 V_low
+ 4.536010000e-07 V_low
+ 4.537000000e-07 V_low
+ 4.537010000e-07 V_low
+ 4.538000000e-07 V_low
+ 4.538010000e-07 V_low
+ 4.539000000e-07 V_low
+ 4.539010000e-07 V_hig
+ 4.540000000e-07 V_hig
+ 4.540010000e-07 V_hig
+ 4.541000000e-07 V_hig
+ 4.541010000e-07 V_hig
+ 4.542000000e-07 V_hig
+ 4.542010000e-07 V_hig
+ 4.543000000e-07 V_hig
+ 4.543010000e-07 V_hig
+ 4.544000000e-07 V_hig
+ 4.544010000e-07 V_hig
+ 4.545000000e-07 V_hig
+ 4.545010000e-07 V_hig
+ 4.546000000e-07 V_hig
+ 4.546010000e-07 V_hig
+ 4.547000000e-07 V_hig
+ 4.547010000e-07 V_hig
+ 4.548000000e-07 V_hig
+ 4.548010000e-07 V_hig
+ 4.549000000e-07 V_hig
+ 4.549010000e-07 V_low
+ 4.550000000e-07 V_low
+ 4.550010000e-07 V_low
+ 4.551000000e-07 V_low
+ 4.551010000e-07 V_low
+ 4.552000000e-07 V_low
+ 4.552010000e-07 V_low
+ 4.553000000e-07 V_low
+ 4.553010000e-07 V_low
+ 4.554000000e-07 V_low
+ 4.554010000e-07 V_low
+ 4.555000000e-07 V_low
+ 4.555010000e-07 V_low
+ 4.556000000e-07 V_low
+ 4.556010000e-07 V_low
+ 4.557000000e-07 V_low
+ 4.557010000e-07 V_low
+ 4.558000000e-07 V_low
+ 4.558010000e-07 V_low
+ 4.559000000e-07 V_low
+ 4.559010000e-07 V_hig
+ 4.560000000e-07 V_hig
+ 4.560010000e-07 V_hig
+ 4.561000000e-07 V_hig
+ 4.561010000e-07 V_hig
+ 4.562000000e-07 V_hig
+ 4.562010000e-07 V_hig
+ 4.563000000e-07 V_hig
+ 4.563010000e-07 V_hig
+ 4.564000000e-07 V_hig
+ 4.564010000e-07 V_hig
+ 4.565000000e-07 V_hig
+ 4.565010000e-07 V_hig
+ 4.566000000e-07 V_hig
+ 4.566010000e-07 V_hig
+ 4.567000000e-07 V_hig
+ 4.567010000e-07 V_hig
+ 4.568000000e-07 V_hig
+ 4.568010000e-07 V_hig
+ 4.569000000e-07 V_hig
+ 4.569010000e-07 V_low
+ 4.570000000e-07 V_low
+ 4.570010000e-07 V_low
+ 4.571000000e-07 V_low
+ 4.571010000e-07 V_low
+ 4.572000000e-07 V_low
+ 4.572010000e-07 V_low
+ 4.573000000e-07 V_low
+ 4.573010000e-07 V_low
+ 4.574000000e-07 V_low
+ 4.574010000e-07 V_low
+ 4.575000000e-07 V_low
+ 4.575010000e-07 V_low
+ 4.576000000e-07 V_low
+ 4.576010000e-07 V_low
+ 4.577000000e-07 V_low
+ 4.577010000e-07 V_low
+ 4.578000000e-07 V_low
+ 4.578010000e-07 V_low
+ 4.579000000e-07 V_low
+ 4.579010000e-07 V_low
+ 4.580000000e-07 V_low
+ 4.580010000e-07 V_low
+ 4.581000000e-07 V_low
+ 4.581010000e-07 V_low
+ 4.582000000e-07 V_low
+ 4.582010000e-07 V_low
+ 4.583000000e-07 V_low
+ 4.583010000e-07 V_low
+ 4.584000000e-07 V_low
+ 4.584010000e-07 V_low
+ 4.585000000e-07 V_low
+ 4.585010000e-07 V_low
+ 4.586000000e-07 V_low
+ 4.586010000e-07 V_low
+ 4.587000000e-07 V_low
+ 4.587010000e-07 V_low
+ 4.588000000e-07 V_low
+ 4.588010000e-07 V_low
+ 4.589000000e-07 V_low
+ 4.589010000e-07 V_low
+ 4.590000000e-07 V_low
+ 4.590010000e-07 V_low
+ 4.591000000e-07 V_low
+ 4.591010000e-07 V_low
+ 4.592000000e-07 V_low
+ 4.592010000e-07 V_low
+ 4.593000000e-07 V_low
+ 4.593010000e-07 V_low
+ 4.594000000e-07 V_low
+ 4.594010000e-07 V_low
+ 4.595000000e-07 V_low
+ 4.595010000e-07 V_low
+ 4.596000000e-07 V_low
+ 4.596010000e-07 V_low
+ 4.597000000e-07 V_low
+ 4.597010000e-07 V_low
+ 4.598000000e-07 V_low
+ 4.598010000e-07 V_low
+ 4.599000000e-07 V_low
+ 4.599010000e-07 V_low
+ 4.600000000e-07 V_low
+ 4.600010000e-07 V_low
+ 4.601000000e-07 V_low
+ 4.601010000e-07 V_low
+ 4.602000000e-07 V_low
+ 4.602010000e-07 V_low
+ 4.603000000e-07 V_low
+ 4.603010000e-07 V_low
+ 4.604000000e-07 V_low
+ 4.604010000e-07 V_low
+ 4.605000000e-07 V_low
+ 4.605010000e-07 V_low
+ 4.606000000e-07 V_low
+ 4.606010000e-07 V_low
+ 4.607000000e-07 V_low
+ 4.607010000e-07 V_low
+ 4.608000000e-07 V_low
+ 4.608010000e-07 V_low
+ 4.609000000e-07 V_low
+ 4.609010000e-07 V_hig
+ 4.610000000e-07 V_hig
+ 4.610010000e-07 V_hig
+ 4.611000000e-07 V_hig
+ 4.611010000e-07 V_hig
+ 4.612000000e-07 V_hig
+ 4.612010000e-07 V_hig
+ 4.613000000e-07 V_hig
+ 4.613010000e-07 V_hig
+ 4.614000000e-07 V_hig
+ 4.614010000e-07 V_hig
+ 4.615000000e-07 V_hig
+ 4.615010000e-07 V_hig
+ 4.616000000e-07 V_hig
+ 4.616010000e-07 V_hig
+ 4.617000000e-07 V_hig
+ 4.617010000e-07 V_hig
+ 4.618000000e-07 V_hig
+ 4.618010000e-07 V_hig
+ 4.619000000e-07 V_hig
+ 4.619010000e-07 V_low
+ 4.620000000e-07 V_low
+ 4.620010000e-07 V_low
+ 4.621000000e-07 V_low
+ 4.621010000e-07 V_low
+ 4.622000000e-07 V_low
+ 4.622010000e-07 V_low
+ 4.623000000e-07 V_low
+ 4.623010000e-07 V_low
+ 4.624000000e-07 V_low
+ 4.624010000e-07 V_low
+ 4.625000000e-07 V_low
+ 4.625010000e-07 V_low
+ 4.626000000e-07 V_low
+ 4.626010000e-07 V_low
+ 4.627000000e-07 V_low
+ 4.627010000e-07 V_low
+ 4.628000000e-07 V_low
+ 4.628010000e-07 V_low
+ 4.629000000e-07 V_low
+ 4.629010000e-07 V_hig
+ 4.630000000e-07 V_hig
+ 4.630010000e-07 V_hig
+ 4.631000000e-07 V_hig
+ 4.631010000e-07 V_hig
+ 4.632000000e-07 V_hig
+ 4.632010000e-07 V_hig
+ 4.633000000e-07 V_hig
+ 4.633010000e-07 V_hig
+ 4.634000000e-07 V_hig
+ 4.634010000e-07 V_hig
+ 4.635000000e-07 V_hig
+ 4.635010000e-07 V_hig
+ 4.636000000e-07 V_hig
+ 4.636010000e-07 V_hig
+ 4.637000000e-07 V_hig
+ 4.637010000e-07 V_hig
+ 4.638000000e-07 V_hig
+ 4.638010000e-07 V_hig
+ 4.639000000e-07 V_hig
+ 4.639010000e-07 V_low
+ 4.640000000e-07 V_low
+ 4.640010000e-07 V_low
+ 4.641000000e-07 V_low
+ 4.641010000e-07 V_low
+ 4.642000000e-07 V_low
+ 4.642010000e-07 V_low
+ 4.643000000e-07 V_low
+ 4.643010000e-07 V_low
+ 4.644000000e-07 V_low
+ 4.644010000e-07 V_low
+ 4.645000000e-07 V_low
+ 4.645010000e-07 V_low
+ 4.646000000e-07 V_low
+ 4.646010000e-07 V_low
+ 4.647000000e-07 V_low
+ 4.647010000e-07 V_low
+ 4.648000000e-07 V_low
+ 4.648010000e-07 V_low
+ 4.649000000e-07 V_low
+ 4.649010000e-07 V_low
+ 4.650000000e-07 V_low
+ 4.650010000e-07 V_low
+ 4.651000000e-07 V_low
+ 4.651010000e-07 V_low
+ 4.652000000e-07 V_low
+ 4.652010000e-07 V_low
+ 4.653000000e-07 V_low
+ 4.653010000e-07 V_low
+ 4.654000000e-07 V_low
+ 4.654010000e-07 V_low
+ 4.655000000e-07 V_low
+ 4.655010000e-07 V_low
+ 4.656000000e-07 V_low
+ 4.656010000e-07 V_low
+ 4.657000000e-07 V_low
+ 4.657010000e-07 V_low
+ 4.658000000e-07 V_low
+ 4.658010000e-07 V_low
+ 4.659000000e-07 V_low
+ 4.659010000e-07 V_low
+ 4.660000000e-07 V_low
+ 4.660010000e-07 V_low
+ 4.661000000e-07 V_low
+ 4.661010000e-07 V_low
+ 4.662000000e-07 V_low
+ 4.662010000e-07 V_low
+ 4.663000000e-07 V_low
+ 4.663010000e-07 V_low
+ 4.664000000e-07 V_low
+ 4.664010000e-07 V_low
+ 4.665000000e-07 V_low
+ 4.665010000e-07 V_low
+ 4.666000000e-07 V_low
+ 4.666010000e-07 V_low
+ 4.667000000e-07 V_low
+ 4.667010000e-07 V_low
+ 4.668000000e-07 V_low
+ 4.668010000e-07 V_low
+ 4.669000000e-07 V_low
+ 4.669010000e-07 V_hig
+ 4.670000000e-07 V_hig
+ 4.670010000e-07 V_hig
+ 4.671000000e-07 V_hig
+ 4.671010000e-07 V_hig
+ 4.672000000e-07 V_hig
+ 4.672010000e-07 V_hig
+ 4.673000000e-07 V_hig
+ 4.673010000e-07 V_hig
+ 4.674000000e-07 V_hig
+ 4.674010000e-07 V_hig
+ 4.675000000e-07 V_hig
+ 4.675010000e-07 V_hig
+ 4.676000000e-07 V_hig
+ 4.676010000e-07 V_hig
+ 4.677000000e-07 V_hig
+ 4.677010000e-07 V_hig
+ 4.678000000e-07 V_hig
+ 4.678010000e-07 V_hig
+ 4.679000000e-07 V_hig
+ 4.679010000e-07 V_hig
+ 4.680000000e-07 V_hig
+ 4.680010000e-07 V_hig
+ 4.681000000e-07 V_hig
+ 4.681010000e-07 V_hig
+ 4.682000000e-07 V_hig
+ 4.682010000e-07 V_hig
+ 4.683000000e-07 V_hig
+ 4.683010000e-07 V_hig
+ 4.684000000e-07 V_hig
+ 4.684010000e-07 V_hig
+ 4.685000000e-07 V_hig
+ 4.685010000e-07 V_hig
+ 4.686000000e-07 V_hig
+ 4.686010000e-07 V_hig
+ 4.687000000e-07 V_hig
+ 4.687010000e-07 V_hig
+ 4.688000000e-07 V_hig
+ 4.688010000e-07 V_hig
+ 4.689000000e-07 V_hig
+ 4.689010000e-07 V_hig
+ 4.690000000e-07 V_hig
+ 4.690010000e-07 V_hig
+ 4.691000000e-07 V_hig
+ 4.691010000e-07 V_hig
+ 4.692000000e-07 V_hig
+ 4.692010000e-07 V_hig
+ 4.693000000e-07 V_hig
+ 4.693010000e-07 V_hig
+ 4.694000000e-07 V_hig
+ 4.694010000e-07 V_hig
+ 4.695000000e-07 V_hig
+ 4.695010000e-07 V_hig
+ 4.696000000e-07 V_hig
+ 4.696010000e-07 V_hig
+ 4.697000000e-07 V_hig
+ 4.697010000e-07 V_hig
+ 4.698000000e-07 V_hig
+ 4.698010000e-07 V_hig
+ 4.699000000e-07 V_hig
+ 4.699010000e-07 V_low
+ 4.700000000e-07 V_low
+ 4.700010000e-07 V_low
+ 4.701000000e-07 V_low
+ 4.701010000e-07 V_low
+ 4.702000000e-07 V_low
+ 4.702010000e-07 V_low
+ 4.703000000e-07 V_low
+ 4.703010000e-07 V_low
+ 4.704000000e-07 V_low
+ 4.704010000e-07 V_low
+ 4.705000000e-07 V_low
+ 4.705010000e-07 V_low
+ 4.706000000e-07 V_low
+ 4.706010000e-07 V_low
+ 4.707000000e-07 V_low
+ 4.707010000e-07 V_low
+ 4.708000000e-07 V_low
+ 4.708010000e-07 V_low
+ 4.709000000e-07 V_low
+ 4.709010000e-07 V_low
+ 4.710000000e-07 V_low
+ 4.710010000e-07 V_low
+ 4.711000000e-07 V_low
+ 4.711010000e-07 V_low
+ 4.712000000e-07 V_low
+ 4.712010000e-07 V_low
+ 4.713000000e-07 V_low
+ 4.713010000e-07 V_low
+ 4.714000000e-07 V_low
+ 4.714010000e-07 V_low
+ 4.715000000e-07 V_low
+ 4.715010000e-07 V_low
+ 4.716000000e-07 V_low
+ 4.716010000e-07 V_low
+ 4.717000000e-07 V_low
+ 4.717010000e-07 V_low
+ 4.718000000e-07 V_low
+ 4.718010000e-07 V_low
+ 4.719000000e-07 V_low
+ 4.719010000e-07 V_hig
+ 4.720000000e-07 V_hig
+ 4.720010000e-07 V_hig
+ 4.721000000e-07 V_hig
+ 4.721010000e-07 V_hig
+ 4.722000000e-07 V_hig
+ 4.722010000e-07 V_hig
+ 4.723000000e-07 V_hig
+ 4.723010000e-07 V_hig
+ 4.724000000e-07 V_hig
+ 4.724010000e-07 V_hig
+ 4.725000000e-07 V_hig
+ 4.725010000e-07 V_hig
+ 4.726000000e-07 V_hig
+ 4.726010000e-07 V_hig
+ 4.727000000e-07 V_hig
+ 4.727010000e-07 V_hig
+ 4.728000000e-07 V_hig
+ 4.728010000e-07 V_hig
+ 4.729000000e-07 V_hig
+ 4.729010000e-07 V_hig
+ 4.730000000e-07 V_hig
+ 4.730010000e-07 V_hig
+ 4.731000000e-07 V_hig
+ 4.731010000e-07 V_hig
+ 4.732000000e-07 V_hig
+ 4.732010000e-07 V_hig
+ 4.733000000e-07 V_hig
+ 4.733010000e-07 V_hig
+ 4.734000000e-07 V_hig
+ 4.734010000e-07 V_hig
+ 4.735000000e-07 V_hig
+ 4.735010000e-07 V_hig
+ 4.736000000e-07 V_hig
+ 4.736010000e-07 V_hig
+ 4.737000000e-07 V_hig
+ 4.737010000e-07 V_hig
+ 4.738000000e-07 V_hig
+ 4.738010000e-07 V_hig
+ 4.739000000e-07 V_hig
+ 4.739010000e-07 V_low
+ 4.740000000e-07 V_low
+ 4.740010000e-07 V_low
+ 4.741000000e-07 V_low
+ 4.741010000e-07 V_low
+ 4.742000000e-07 V_low
+ 4.742010000e-07 V_low
+ 4.743000000e-07 V_low
+ 4.743010000e-07 V_low
+ 4.744000000e-07 V_low
+ 4.744010000e-07 V_low
+ 4.745000000e-07 V_low
+ 4.745010000e-07 V_low
+ 4.746000000e-07 V_low
+ 4.746010000e-07 V_low
+ 4.747000000e-07 V_low
+ 4.747010000e-07 V_low
+ 4.748000000e-07 V_low
+ 4.748010000e-07 V_low
+ 4.749000000e-07 V_low
+ 4.749010000e-07 V_low
+ 4.750000000e-07 V_low
+ 4.750010000e-07 V_low
+ 4.751000000e-07 V_low
+ 4.751010000e-07 V_low
+ 4.752000000e-07 V_low
+ 4.752010000e-07 V_low
+ 4.753000000e-07 V_low
+ 4.753010000e-07 V_low
+ 4.754000000e-07 V_low
+ 4.754010000e-07 V_low
+ 4.755000000e-07 V_low
+ 4.755010000e-07 V_low
+ 4.756000000e-07 V_low
+ 4.756010000e-07 V_low
+ 4.757000000e-07 V_low
+ 4.757010000e-07 V_low
+ 4.758000000e-07 V_low
+ 4.758010000e-07 V_low
+ 4.759000000e-07 V_low
+ 4.759010000e-07 V_low
+ 4.760000000e-07 V_low
+ 4.760010000e-07 V_low
+ 4.761000000e-07 V_low
+ 4.761010000e-07 V_low
+ 4.762000000e-07 V_low
+ 4.762010000e-07 V_low
+ 4.763000000e-07 V_low
+ 4.763010000e-07 V_low
+ 4.764000000e-07 V_low
+ 4.764010000e-07 V_low
+ 4.765000000e-07 V_low
+ 4.765010000e-07 V_low
+ 4.766000000e-07 V_low
+ 4.766010000e-07 V_low
+ 4.767000000e-07 V_low
+ 4.767010000e-07 V_low
+ 4.768000000e-07 V_low
+ 4.768010000e-07 V_low
+ 4.769000000e-07 V_low
+ 4.769010000e-07 V_hig
+ 4.770000000e-07 V_hig
+ 4.770010000e-07 V_hig
+ 4.771000000e-07 V_hig
+ 4.771010000e-07 V_hig
+ 4.772000000e-07 V_hig
+ 4.772010000e-07 V_hig
+ 4.773000000e-07 V_hig
+ 4.773010000e-07 V_hig
+ 4.774000000e-07 V_hig
+ 4.774010000e-07 V_hig
+ 4.775000000e-07 V_hig
+ 4.775010000e-07 V_hig
+ 4.776000000e-07 V_hig
+ 4.776010000e-07 V_hig
+ 4.777000000e-07 V_hig
+ 4.777010000e-07 V_hig
+ 4.778000000e-07 V_hig
+ 4.778010000e-07 V_hig
+ 4.779000000e-07 V_hig
+ 4.779010000e-07 V_hig
+ 4.780000000e-07 V_hig
+ 4.780010000e-07 V_hig
+ 4.781000000e-07 V_hig
+ 4.781010000e-07 V_hig
+ 4.782000000e-07 V_hig
+ 4.782010000e-07 V_hig
+ 4.783000000e-07 V_hig
+ 4.783010000e-07 V_hig
+ 4.784000000e-07 V_hig
+ 4.784010000e-07 V_hig
+ 4.785000000e-07 V_hig
+ 4.785010000e-07 V_hig
+ 4.786000000e-07 V_hig
+ 4.786010000e-07 V_hig
+ 4.787000000e-07 V_hig
+ 4.787010000e-07 V_hig
+ 4.788000000e-07 V_hig
+ 4.788010000e-07 V_hig
+ 4.789000000e-07 V_hig
+ 4.789010000e-07 V_hig
+ 4.790000000e-07 V_hig
+ 4.790010000e-07 V_hig
+ 4.791000000e-07 V_hig
+ 4.791010000e-07 V_hig
+ 4.792000000e-07 V_hig
+ 4.792010000e-07 V_hig
+ 4.793000000e-07 V_hig
+ 4.793010000e-07 V_hig
+ 4.794000000e-07 V_hig
+ 4.794010000e-07 V_hig
+ 4.795000000e-07 V_hig
+ 4.795010000e-07 V_hig
+ 4.796000000e-07 V_hig
+ 4.796010000e-07 V_hig
+ 4.797000000e-07 V_hig
+ 4.797010000e-07 V_hig
+ 4.798000000e-07 V_hig
+ 4.798010000e-07 V_hig
+ 4.799000000e-07 V_hig
+ 4.799010000e-07 V_hig
+ 4.800000000e-07 V_hig
+ 4.800010000e-07 V_hig
+ 4.801000000e-07 V_hig
+ 4.801010000e-07 V_hig
+ 4.802000000e-07 V_hig
+ 4.802010000e-07 V_hig
+ 4.803000000e-07 V_hig
+ 4.803010000e-07 V_hig
+ 4.804000000e-07 V_hig
+ 4.804010000e-07 V_hig
+ 4.805000000e-07 V_hig
+ 4.805010000e-07 V_hig
+ 4.806000000e-07 V_hig
+ 4.806010000e-07 V_hig
+ 4.807000000e-07 V_hig
+ 4.807010000e-07 V_hig
+ 4.808000000e-07 V_hig
+ 4.808010000e-07 V_hig
+ 4.809000000e-07 V_hig
+ 4.809010000e-07 V_low
+ 4.810000000e-07 V_low
+ 4.810010000e-07 V_low
+ 4.811000000e-07 V_low
+ 4.811010000e-07 V_low
+ 4.812000000e-07 V_low
+ 4.812010000e-07 V_low
+ 4.813000000e-07 V_low
+ 4.813010000e-07 V_low
+ 4.814000000e-07 V_low
+ 4.814010000e-07 V_low
+ 4.815000000e-07 V_low
+ 4.815010000e-07 V_low
+ 4.816000000e-07 V_low
+ 4.816010000e-07 V_low
+ 4.817000000e-07 V_low
+ 4.817010000e-07 V_low
+ 4.818000000e-07 V_low
+ 4.818010000e-07 V_low
+ 4.819000000e-07 V_low
+ 4.819010000e-07 V_low
+ 4.820000000e-07 V_low
+ 4.820010000e-07 V_low
+ 4.821000000e-07 V_low
+ 4.821010000e-07 V_low
+ 4.822000000e-07 V_low
+ 4.822010000e-07 V_low
+ 4.823000000e-07 V_low
+ 4.823010000e-07 V_low
+ 4.824000000e-07 V_low
+ 4.824010000e-07 V_low
+ 4.825000000e-07 V_low
+ 4.825010000e-07 V_low
+ 4.826000000e-07 V_low
+ 4.826010000e-07 V_low
+ 4.827000000e-07 V_low
+ 4.827010000e-07 V_low
+ 4.828000000e-07 V_low
+ 4.828010000e-07 V_low
+ 4.829000000e-07 V_low
+ 4.829010000e-07 V_hig
+ 4.830000000e-07 V_hig
+ 4.830010000e-07 V_hig
+ 4.831000000e-07 V_hig
+ 4.831010000e-07 V_hig
+ 4.832000000e-07 V_hig
+ 4.832010000e-07 V_hig
+ 4.833000000e-07 V_hig
+ 4.833010000e-07 V_hig
+ 4.834000000e-07 V_hig
+ 4.834010000e-07 V_hig
+ 4.835000000e-07 V_hig
+ 4.835010000e-07 V_hig
+ 4.836000000e-07 V_hig
+ 4.836010000e-07 V_hig
+ 4.837000000e-07 V_hig
+ 4.837010000e-07 V_hig
+ 4.838000000e-07 V_hig
+ 4.838010000e-07 V_hig
+ 4.839000000e-07 V_hig
+ 4.839010000e-07 V_hig
+ 4.840000000e-07 V_hig
+ 4.840010000e-07 V_hig
+ 4.841000000e-07 V_hig
+ 4.841010000e-07 V_hig
+ 4.842000000e-07 V_hig
+ 4.842010000e-07 V_hig
+ 4.843000000e-07 V_hig
+ 4.843010000e-07 V_hig
+ 4.844000000e-07 V_hig
+ 4.844010000e-07 V_hig
+ 4.845000000e-07 V_hig
+ 4.845010000e-07 V_hig
+ 4.846000000e-07 V_hig
+ 4.846010000e-07 V_hig
+ 4.847000000e-07 V_hig
+ 4.847010000e-07 V_hig
+ 4.848000000e-07 V_hig
+ 4.848010000e-07 V_hig
+ 4.849000000e-07 V_hig
+ 4.849010000e-07 V_low
+ 4.850000000e-07 V_low
+ 4.850010000e-07 V_low
+ 4.851000000e-07 V_low
+ 4.851010000e-07 V_low
+ 4.852000000e-07 V_low
+ 4.852010000e-07 V_low
+ 4.853000000e-07 V_low
+ 4.853010000e-07 V_low
+ 4.854000000e-07 V_low
+ 4.854010000e-07 V_low
+ 4.855000000e-07 V_low
+ 4.855010000e-07 V_low
+ 4.856000000e-07 V_low
+ 4.856010000e-07 V_low
+ 4.857000000e-07 V_low
+ 4.857010000e-07 V_low
+ 4.858000000e-07 V_low
+ 4.858010000e-07 V_low
+ 4.859000000e-07 V_low
+ 4.859010000e-07 V_hig
+ 4.860000000e-07 V_hig
+ 4.860010000e-07 V_hig
+ 4.861000000e-07 V_hig
+ 4.861010000e-07 V_hig
+ 4.862000000e-07 V_hig
+ 4.862010000e-07 V_hig
+ 4.863000000e-07 V_hig
+ 4.863010000e-07 V_hig
+ 4.864000000e-07 V_hig
+ 4.864010000e-07 V_hig
+ 4.865000000e-07 V_hig
+ 4.865010000e-07 V_hig
+ 4.866000000e-07 V_hig
+ 4.866010000e-07 V_hig
+ 4.867000000e-07 V_hig
+ 4.867010000e-07 V_hig
+ 4.868000000e-07 V_hig
+ 4.868010000e-07 V_hig
+ 4.869000000e-07 V_hig
+ 4.869010000e-07 V_hig
+ 4.870000000e-07 V_hig
+ 4.870010000e-07 V_hig
+ 4.871000000e-07 V_hig
+ 4.871010000e-07 V_hig
+ 4.872000000e-07 V_hig
+ 4.872010000e-07 V_hig
+ 4.873000000e-07 V_hig
+ 4.873010000e-07 V_hig
+ 4.874000000e-07 V_hig
+ 4.874010000e-07 V_hig
+ 4.875000000e-07 V_hig
+ 4.875010000e-07 V_hig
+ 4.876000000e-07 V_hig
+ 4.876010000e-07 V_hig
+ 4.877000000e-07 V_hig
+ 4.877010000e-07 V_hig
+ 4.878000000e-07 V_hig
+ 4.878010000e-07 V_hig
+ 4.879000000e-07 V_hig
+ 4.879010000e-07 V_low
+ 4.880000000e-07 V_low
+ 4.880010000e-07 V_low
+ 4.881000000e-07 V_low
+ 4.881010000e-07 V_low
+ 4.882000000e-07 V_low
+ 4.882010000e-07 V_low
+ 4.883000000e-07 V_low
+ 4.883010000e-07 V_low
+ 4.884000000e-07 V_low
+ 4.884010000e-07 V_low
+ 4.885000000e-07 V_low
+ 4.885010000e-07 V_low
+ 4.886000000e-07 V_low
+ 4.886010000e-07 V_low
+ 4.887000000e-07 V_low
+ 4.887010000e-07 V_low
+ 4.888000000e-07 V_low
+ 4.888010000e-07 V_low
+ 4.889000000e-07 V_low
+ 4.889010000e-07 V_low
+ 4.890000000e-07 V_low
+ 4.890010000e-07 V_low
+ 4.891000000e-07 V_low
+ 4.891010000e-07 V_low
+ 4.892000000e-07 V_low
+ 4.892010000e-07 V_low
+ 4.893000000e-07 V_low
+ 4.893010000e-07 V_low
+ 4.894000000e-07 V_low
+ 4.894010000e-07 V_low
+ 4.895000000e-07 V_low
+ 4.895010000e-07 V_low
+ 4.896000000e-07 V_low
+ 4.896010000e-07 V_low
+ 4.897000000e-07 V_low
+ 4.897010000e-07 V_low
+ 4.898000000e-07 V_low
+ 4.898010000e-07 V_low
+ 4.899000000e-07 V_low
+ 4.899010000e-07 V_low
+ 4.900000000e-07 V_low
+ 4.900010000e-07 V_low
+ 4.901000000e-07 V_low
+ 4.901010000e-07 V_low
+ 4.902000000e-07 V_low
+ 4.902010000e-07 V_low
+ 4.903000000e-07 V_low
+ 4.903010000e-07 V_low
+ 4.904000000e-07 V_low
+ 4.904010000e-07 V_low
+ 4.905000000e-07 V_low
+ 4.905010000e-07 V_low
+ 4.906000000e-07 V_low
+ 4.906010000e-07 V_low
+ 4.907000000e-07 V_low
+ 4.907010000e-07 V_low
+ 4.908000000e-07 V_low
+ 4.908010000e-07 V_low
+ 4.909000000e-07 V_low
+ 4.909010000e-07 V_hig
+ 4.910000000e-07 V_hig
+ 4.910010000e-07 V_hig
+ 4.911000000e-07 V_hig
+ 4.911010000e-07 V_hig
+ 4.912000000e-07 V_hig
+ 4.912010000e-07 V_hig
+ 4.913000000e-07 V_hig
+ 4.913010000e-07 V_hig
+ 4.914000000e-07 V_hig
+ 4.914010000e-07 V_hig
+ 4.915000000e-07 V_hig
+ 4.915010000e-07 V_hig
+ 4.916000000e-07 V_hig
+ 4.916010000e-07 V_hig
+ 4.917000000e-07 V_hig
+ 4.917010000e-07 V_hig
+ 4.918000000e-07 V_hig
+ 4.918010000e-07 V_hig
+ 4.919000000e-07 V_hig
+ 4.919010000e-07 V_low
+ 4.920000000e-07 V_low
+ 4.920010000e-07 V_low
+ 4.921000000e-07 V_low
+ 4.921010000e-07 V_low
+ 4.922000000e-07 V_low
+ 4.922010000e-07 V_low
+ 4.923000000e-07 V_low
+ 4.923010000e-07 V_low
+ 4.924000000e-07 V_low
+ 4.924010000e-07 V_low
+ 4.925000000e-07 V_low
+ 4.925010000e-07 V_low
+ 4.926000000e-07 V_low
+ 4.926010000e-07 V_low
+ 4.927000000e-07 V_low
+ 4.927010000e-07 V_low
+ 4.928000000e-07 V_low
+ 4.928010000e-07 V_low
+ 4.929000000e-07 V_low
+ 4.929010000e-07 V_low
+ 4.930000000e-07 V_low
+ 4.930010000e-07 V_low
+ 4.931000000e-07 V_low
+ 4.931010000e-07 V_low
+ 4.932000000e-07 V_low
+ 4.932010000e-07 V_low
+ 4.933000000e-07 V_low
+ 4.933010000e-07 V_low
+ 4.934000000e-07 V_low
+ 4.934010000e-07 V_low
+ 4.935000000e-07 V_low
+ 4.935010000e-07 V_low
+ 4.936000000e-07 V_low
+ 4.936010000e-07 V_low
+ 4.937000000e-07 V_low
+ 4.937010000e-07 V_low
+ 4.938000000e-07 V_low
+ 4.938010000e-07 V_low
+ 4.939000000e-07 V_low
+ 4.939010000e-07 V_low
+ 4.940000000e-07 V_low
+ 4.940010000e-07 V_low
+ 4.941000000e-07 V_low
+ 4.941010000e-07 V_low
+ 4.942000000e-07 V_low
+ 4.942010000e-07 V_low
+ 4.943000000e-07 V_low
+ 4.943010000e-07 V_low
+ 4.944000000e-07 V_low
+ 4.944010000e-07 V_low
+ 4.945000000e-07 V_low
+ 4.945010000e-07 V_low
+ 4.946000000e-07 V_low
+ 4.946010000e-07 V_low
+ 4.947000000e-07 V_low
+ 4.947010000e-07 V_low
+ 4.948000000e-07 V_low
+ 4.948010000e-07 V_low
+ 4.949000000e-07 V_low
+ 4.949010000e-07 V_hig
+ 4.950000000e-07 V_hig
+ 4.950010000e-07 V_hig
+ 4.951000000e-07 V_hig
+ 4.951010000e-07 V_hig
+ 4.952000000e-07 V_hig
+ 4.952010000e-07 V_hig
+ 4.953000000e-07 V_hig
+ 4.953010000e-07 V_hig
+ 4.954000000e-07 V_hig
+ 4.954010000e-07 V_hig
+ 4.955000000e-07 V_hig
+ 4.955010000e-07 V_hig
+ 4.956000000e-07 V_hig
+ 4.956010000e-07 V_hig
+ 4.957000000e-07 V_hig
+ 4.957010000e-07 V_hig
+ 4.958000000e-07 V_hig
+ 4.958010000e-07 V_hig
+ 4.959000000e-07 V_hig
+ 4.959010000e-07 V_hig
+ 4.960000000e-07 V_hig
+ 4.960010000e-07 V_hig
+ 4.961000000e-07 V_hig
+ 4.961010000e-07 V_hig
+ 4.962000000e-07 V_hig
+ 4.962010000e-07 V_hig
+ 4.963000000e-07 V_hig
+ 4.963010000e-07 V_hig
+ 4.964000000e-07 V_hig
+ 4.964010000e-07 V_hig
+ 4.965000000e-07 V_hig
+ 4.965010000e-07 V_hig
+ 4.966000000e-07 V_hig
+ 4.966010000e-07 V_hig
+ 4.967000000e-07 V_hig
+ 4.967010000e-07 V_hig
+ 4.968000000e-07 V_hig
+ 4.968010000e-07 V_hig
+ 4.969000000e-07 V_hig
+ 4.969010000e-07 V_hig
+ 4.970000000e-07 V_hig
+ 4.970010000e-07 V_hig
+ 4.971000000e-07 V_hig
+ 4.971010000e-07 V_hig
+ 4.972000000e-07 V_hig
+ 4.972010000e-07 V_hig
+ 4.973000000e-07 V_hig
+ 4.973010000e-07 V_hig
+ 4.974000000e-07 V_hig
+ 4.974010000e-07 V_hig
+ 4.975000000e-07 V_hig
+ 4.975010000e-07 V_hig
+ 4.976000000e-07 V_hig
+ 4.976010000e-07 V_hig
+ 4.977000000e-07 V_hig
+ 4.977010000e-07 V_hig
+ 4.978000000e-07 V_hig
+ 4.978010000e-07 V_hig
+ 4.979000000e-07 V_hig
+ 4.979010000e-07 V_hig
+ 4.980000000e-07 V_hig
+ 4.980010000e-07 V_hig
+ 4.981000000e-07 V_hig
+ 4.981010000e-07 V_hig
+ 4.982000000e-07 V_hig
+ 4.982010000e-07 V_hig
+ 4.983000000e-07 V_hig
+ 4.983010000e-07 V_hig
+ 4.984000000e-07 V_hig
+ 4.984010000e-07 V_hig
+ 4.985000000e-07 V_hig
+ 4.985010000e-07 V_hig
+ 4.986000000e-07 V_hig
+ 4.986010000e-07 V_hig
+ 4.987000000e-07 V_hig
+ 4.987010000e-07 V_hig
+ 4.988000000e-07 V_hig
+ 4.988010000e-07 V_hig
+ 4.989000000e-07 V_hig
+ 4.989010000e-07 V_low
+ 4.990000000e-07 V_low
+ 4.990010000e-07 V_low
+ 4.991000000e-07 V_low
+ 4.991010000e-07 V_low
+ 4.992000000e-07 V_low
+ 4.992010000e-07 V_low
+ 4.993000000e-07 V_low
+ 4.993010000e-07 V_low
+ 4.994000000e-07 V_low
+ 4.994010000e-07 V_low
+ 4.995000000e-07 V_low
+ 4.995010000e-07 V_low
+ 4.996000000e-07 V_low
+ 4.996010000e-07 V_low
+ 4.997000000e-07 V_low
+ 4.997010000e-07 V_low
+ 4.998000000e-07 V_low
+ 4.998010000e-07 V_low
+ 4.999000000e-07 V_low
+ 4.999010000e-07 V_hig
+ 5.000000000e-07 V_hig
+ 5.000010000e-07 V_hig
+ 5.001000000e-07 V_hig
+ 5.001010000e-07 V_hig
+ 5.002000000e-07 V_hig
+ 5.002010000e-07 V_hig
+ 5.003000000e-07 V_hig
+ 5.003010000e-07 V_hig
+ 5.004000000e-07 V_hig
+ 5.004010000e-07 V_hig
+ 5.005000000e-07 V_hig
+ 5.005010000e-07 V_hig
+ 5.006000000e-07 V_hig
+ 5.006010000e-07 V_hig
+ 5.007000000e-07 V_hig
+ 5.007010000e-07 V_hig
+ 5.008000000e-07 V_hig
+ 5.008010000e-07 V_hig
+ 5.009000000e-07 V_hig
+ 5.009010000e-07 V_low
+ 5.010000000e-07 V_low
+ 5.010010000e-07 V_low
+ 5.011000000e-07 V_low
+ 5.011010000e-07 V_low
+ 5.012000000e-07 V_low
+ 5.012010000e-07 V_low
+ 5.013000000e-07 V_low
+ 5.013010000e-07 V_low
+ 5.014000000e-07 V_low
+ 5.014010000e-07 V_low
+ 5.015000000e-07 V_low
+ 5.015010000e-07 V_low
+ 5.016000000e-07 V_low
+ 5.016010000e-07 V_low
+ 5.017000000e-07 V_low
+ 5.017010000e-07 V_low
+ 5.018000000e-07 V_low
+ 5.018010000e-07 V_low
+ 5.019000000e-07 V_low
+ 5.019010000e-07 V_hig
+ 5.020000000e-07 V_hig
+ 5.020010000e-07 V_hig
+ 5.021000000e-07 V_hig
+ 5.021010000e-07 V_hig
+ 5.022000000e-07 V_hig
+ 5.022010000e-07 V_hig
+ 5.023000000e-07 V_hig
+ 5.023010000e-07 V_hig
+ 5.024000000e-07 V_hig
+ 5.024010000e-07 V_hig
+ 5.025000000e-07 V_hig
+ 5.025010000e-07 V_hig
+ 5.026000000e-07 V_hig
+ 5.026010000e-07 V_hig
+ 5.027000000e-07 V_hig
+ 5.027010000e-07 V_hig
+ 5.028000000e-07 V_hig
+ 5.028010000e-07 V_hig
+ 5.029000000e-07 V_hig
+ 5.029010000e-07 V_low
+ 5.030000000e-07 V_low
+ 5.030010000e-07 V_low
+ 5.031000000e-07 V_low
+ 5.031010000e-07 V_low
+ 5.032000000e-07 V_low
+ 5.032010000e-07 V_low
+ 5.033000000e-07 V_low
+ 5.033010000e-07 V_low
+ 5.034000000e-07 V_low
+ 5.034010000e-07 V_low
+ 5.035000000e-07 V_low
+ 5.035010000e-07 V_low
+ 5.036000000e-07 V_low
+ 5.036010000e-07 V_low
+ 5.037000000e-07 V_low
+ 5.037010000e-07 V_low
+ 5.038000000e-07 V_low
+ 5.038010000e-07 V_low
+ 5.039000000e-07 V_low
+ 5.039010000e-07 V_hig
+ 5.040000000e-07 V_hig
+ 5.040010000e-07 V_hig
+ 5.041000000e-07 V_hig
+ 5.041010000e-07 V_hig
+ 5.042000000e-07 V_hig
+ 5.042010000e-07 V_hig
+ 5.043000000e-07 V_hig
+ 5.043010000e-07 V_hig
+ 5.044000000e-07 V_hig
+ 5.044010000e-07 V_hig
+ 5.045000000e-07 V_hig
+ 5.045010000e-07 V_hig
+ 5.046000000e-07 V_hig
+ 5.046010000e-07 V_hig
+ 5.047000000e-07 V_hig
+ 5.047010000e-07 V_hig
+ 5.048000000e-07 V_hig
+ 5.048010000e-07 V_hig
+ 5.049000000e-07 V_hig
+ 5.049010000e-07 V_hig
+ 5.050000000e-07 V_hig
+ 5.050010000e-07 V_hig
+ 5.051000000e-07 V_hig
+ 5.051010000e-07 V_hig
+ 5.052000000e-07 V_hig
+ 5.052010000e-07 V_hig
+ 5.053000000e-07 V_hig
+ 5.053010000e-07 V_hig
+ 5.054000000e-07 V_hig
+ 5.054010000e-07 V_hig
+ 5.055000000e-07 V_hig
+ 5.055010000e-07 V_hig
+ 5.056000000e-07 V_hig
+ 5.056010000e-07 V_hig
+ 5.057000000e-07 V_hig
+ 5.057010000e-07 V_hig
+ 5.058000000e-07 V_hig
+ 5.058010000e-07 V_hig
+ 5.059000000e-07 V_hig
+ 5.059010000e-07 V_hig
+ 5.060000000e-07 V_hig
+ 5.060010000e-07 V_hig
+ 5.061000000e-07 V_hig
+ 5.061010000e-07 V_hig
+ 5.062000000e-07 V_hig
+ 5.062010000e-07 V_hig
+ 5.063000000e-07 V_hig
+ 5.063010000e-07 V_hig
+ 5.064000000e-07 V_hig
+ 5.064010000e-07 V_hig
+ 5.065000000e-07 V_hig
+ 5.065010000e-07 V_hig
+ 5.066000000e-07 V_hig
+ 5.066010000e-07 V_hig
+ 5.067000000e-07 V_hig
+ 5.067010000e-07 V_hig
+ 5.068000000e-07 V_hig
+ 5.068010000e-07 V_hig
+ 5.069000000e-07 V_hig
+ 5.069010000e-07 V_hig
+ 5.070000000e-07 V_hig
+ 5.070010000e-07 V_hig
+ 5.071000000e-07 V_hig
+ 5.071010000e-07 V_hig
+ 5.072000000e-07 V_hig
+ 5.072010000e-07 V_hig
+ 5.073000000e-07 V_hig
+ 5.073010000e-07 V_hig
+ 5.074000000e-07 V_hig
+ 5.074010000e-07 V_hig
+ 5.075000000e-07 V_hig
+ 5.075010000e-07 V_hig
+ 5.076000000e-07 V_hig
+ 5.076010000e-07 V_hig
+ 5.077000000e-07 V_hig
+ 5.077010000e-07 V_hig
+ 5.078000000e-07 V_hig
+ 5.078010000e-07 V_hig
+ 5.079000000e-07 V_hig
+ 5.079010000e-07 V_hig
+ 5.080000000e-07 V_hig
+ 5.080010000e-07 V_hig
+ 5.081000000e-07 V_hig
+ 5.081010000e-07 V_hig
+ 5.082000000e-07 V_hig
+ 5.082010000e-07 V_hig
+ 5.083000000e-07 V_hig
+ 5.083010000e-07 V_hig
+ 5.084000000e-07 V_hig
+ 5.084010000e-07 V_hig
+ 5.085000000e-07 V_hig
+ 5.085010000e-07 V_hig
+ 5.086000000e-07 V_hig
+ 5.086010000e-07 V_hig
+ 5.087000000e-07 V_hig
+ 5.087010000e-07 V_hig
+ 5.088000000e-07 V_hig
+ 5.088010000e-07 V_hig
+ 5.089000000e-07 V_hig
+ 5.089010000e-07 V_low
+ 5.090000000e-07 V_low
+ 5.090010000e-07 V_low
+ 5.091000000e-07 V_low
+ 5.091010000e-07 V_low
+ 5.092000000e-07 V_low
+ 5.092010000e-07 V_low
+ 5.093000000e-07 V_low
+ 5.093010000e-07 V_low
+ 5.094000000e-07 V_low
+ 5.094010000e-07 V_low
+ 5.095000000e-07 V_low
+ 5.095010000e-07 V_low
+ 5.096000000e-07 V_low
+ 5.096010000e-07 V_low
+ 5.097000000e-07 V_low
+ 5.097010000e-07 V_low
+ 5.098000000e-07 V_low
+ 5.098010000e-07 V_low
+ 5.099000000e-07 V_low
+ 5.099010000e-07 V_hig
+ 5.100000000e-07 V_hig
+ 5.100010000e-07 V_hig
+ 5.101000000e-07 V_hig
+ 5.101010000e-07 V_hig
+ 5.102000000e-07 V_hig
+ 5.102010000e-07 V_hig
+ 5.103000000e-07 V_hig
+ 5.103010000e-07 V_hig
+ 5.104000000e-07 V_hig
+ 5.104010000e-07 V_hig
+ 5.105000000e-07 V_hig
+ 5.105010000e-07 V_hig
+ 5.106000000e-07 V_hig
+ 5.106010000e-07 V_hig
+ 5.107000000e-07 V_hig
+ 5.107010000e-07 V_hig
+ 5.108000000e-07 V_hig
+ 5.108010000e-07 V_hig
+ 5.109000000e-07 V_hig
+ 5.109010000e-07 V_hig
+ 5.110000000e-07 V_hig
+ 5.110010000e-07 V_hig
+ 5.111000000e-07 V_hig
+ 5.111010000e-07 V_hig
+ 5.112000000e-07 V_hig
+ 5.112010000e-07 V_hig
+ 5.113000000e-07 V_hig
+ 5.113010000e-07 V_hig
+ 5.114000000e-07 V_hig
+ 5.114010000e-07 V_hig
+ 5.115000000e-07 V_hig
+ 5.115010000e-07 V_hig
+ 5.116000000e-07 V_hig
+ 5.116010000e-07 V_hig
+ 5.117000000e-07 V_hig
+ 5.117010000e-07 V_hig
+ 5.118000000e-07 V_hig
+ 5.118010000e-07 V_hig
+ 5.119000000e-07 V_hig
+ 5.119010000e-07 V_hig
+ 5.120000000e-07 V_hig
+ 5.120010000e-07 V_hig
+ 5.121000000e-07 V_hig
+ 5.121010000e-07 V_hig
+ 5.122000000e-07 V_hig
+ 5.122010000e-07 V_hig
+ 5.123000000e-07 V_hig
+ 5.123010000e-07 V_hig
+ 5.124000000e-07 V_hig
+ 5.124010000e-07 V_hig
+ 5.125000000e-07 V_hig
+ 5.125010000e-07 V_hig
+ 5.126000000e-07 V_hig
+ 5.126010000e-07 V_hig
+ 5.127000000e-07 V_hig
+ 5.127010000e-07 V_hig
+ 5.128000000e-07 V_hig
+ 5.128010000e-07 V_hig
+ 5.129000000e-07 V_hig
+ 5.129010000e-07 V_low
+ 5.130000000e-07 V_low
+ 5.130010000e-07 V_low
+ 5.131000000e-07 V_low
+ 5.131010000e-07 V_low
+ 5.132000000e-07 V_low
+ 5.132010000e-07 V_low
+ 5.133000000e-07 V_low
+ 5.133010000e-07 V_low
+ 5.134000000e-07 V_low
+ 5.134010000e-07 V_low
+ 5.135000000e-07 V_low
+ 5.135010000e-07 V_low
+ 5.136000000e-07 V_low
+ 5.136010000e-07 V_low
+ 5.137000000e-07 V_low
+ 5.137010000e-07 V_low
+ 5.138000000e-07 V_low
+ 5.138010000e-07 V_low
+ 5.139000000e-07 V_low
+ 5.139010000e-07 V_hig
+ 5.140000000e-07 V_hig
+ 5.140010000e-07 V_hig
+ 5.141000000e-07 V_hig
+ 5.141010000e-07 V_hig
+ 5.142000000e-07 V_hig
+ 5.142010000e-07 V_hig
+ 5.143000000e-07 V_hig
+ 5.143010000e-07 V_hig
+ 5.144000000e-07 V_hig
+ 5.144010000e-07 V_hig
+ 5.145000000e-07 V_hig
+ 5.145010000e-07 V_hig
+ 5.146000000e-07 V_hig
+ 5.146010000e-07 V_hig
+ 5.147000000e-07 V_hig
+ 5.147010000e-07 V_hig
+ 5.148000000e-07 V_hig
+ 5.148010000e-07 V_hig
+ 5.149000000e-07 V_hig
+ 5.149010000e-07 V_hig
+ 5.150000000e-07 V_hig
+ 5.150010000e-07 V_hig
+ 5.151000000e-07 V_hig
+ 5.151010000e-07 V_hig
+ 5.152000000e-07 V_hig
+ 5.152010000e-07 V_hig
+ 5.153000000e-07 V_hig
+ 5.153010000e-07 V_hig
+ 5.154000000e-07 V_hig
+ 5.154010000e-07 V_hig
+ 5.155000000e-07 V_hig
+ 5.155010000e-07 V_hig
+ 5.156000000e-07 V_hig
+ 5.156010000e-07 V_hig
+ 5.157000000e-07 V_hig
+ 5.157010000e-07 V_hig
+ 5.158000000e-07 V_hig
+ 5.158010000e-07 V_hig
+ 5.159000000e-07 V_hig
+ 5.159010000e-07 V_low
+ 5.160000000e-07 V_low
+ 5.160010000e-07 V_low
+ 5.161000000e-07 V_low
+ 5.161010000e-07 V_low
+ 5.162000000e-07 V_low
+ 5.162010000e-07 V_low
+ 5.163000000e-07 V_low
+ 5.163010000e-07 V_low
+ 5.164000000e-07 V_low
+ 5.164010000e-07 V_low
+ 5.165000000e-07 V_low
+ 5.165010000e-07 V_low
+ 5.166000000e-07 V_low
+ 5.166010000e-07 V_low
+ 5.167000000e-07 V_low
+ 5.167010000e-07 V_low
+ 5.168000000e-07 V_low
+ 5.168010000e-07 V_low
+ 5.169000000e-07 V_low
+ 5.169010000e-07 V_hig
+ 5.170000000e-07 V_hig
+ 5.170010000e-07 V_hig
+ 5.171000000e-07 V_hig
+ 5.171010000e-07 V_hig
+ 5.172000000e-07 V_hig
+ 5.172010000e-07 V_hig
+ 5.173000000e-07 V_hig
+ 5.173010000e-07 V_hig
+ 5.174000000e-07 V_hig
+ 5.174010000e-07 V_hig
+ 5.175000000e-07 V_hig
+ 5.175010000e-07 V_hig
+ 5.176000000e-07 V_hig
+ 5.176010000e-07 V_hig
+ 5.177000000e-07 V_hig
+ 5.177010000e-07 V_hig
+ 5.178000000e-07 V_hig
+ 5.178010000e-07 V_hig
+ 5.179000000e-07 V_hig
+ 5.179010000e-07 V_hig
+ 5.180000000e-07 V_hig
+ 5.180010000e-07 V_hig
+ 5.181000000e-07 V_hig
+ 5.181010000e-07 V_hig
+ 5.182000000e-07 V_hig
+ 5.182010000e-07 V_hig
+ 5.183000000e-07 V_hig
+ 5.183010000e-07 V_hig
+ 5.184000000e-07 V_hig
+ 5.184010000e-07 V_hig
+ 5.185000000e-07 V_hig
+ 5.185010000e-07 V_hig
+ 5.186000000e-07 V_hig
+ 5.186010000e-07 V_hig
+ 5.187000000e-07 V_hig
+ 5.187010000e-07 V_hig
+ 5.188000000e-07 V_hig
+ 5.188010000e-07 V_hig
+ 5.189000000e-07 V_hig
+ 5.189010000e-07 V_hig
+ 5.190000000e-07 V_hig
+ 5.190010000e-07 V_hig
+ 5.191000000e-07 V_hig
+ 5.191010000e-07 V_hig
+ 5.192000000e-07 V_hig
+ 5.192010000e-07 V_hig
+ 5.193000000e-07 V_hig
+ 5.193010000e-07 V_hig
+ 5.194000000e-07 V_hig
+ 5.194010000e-07 V_hig
+ 5.195000000e-07 V_hig
+ 5.195010000e-07 V_hig
+ 5.196000000e-07 V_hig
+ 5.196010000e-07 V_hig
+ 5.197000000e-07 V_hig
+ 5.197010000e-07 V_hig
+ 5.198000000e-07 V_hig
+ 5.198010000e-07 V_hig
+ 5.199000000e-07 V_hig
+ 5.199010000e-07 V_hig
+ 5.200000000e-07 V_hig
+ 5.200010000e-07 V_hig
+ 5.201000000e-07 V_hig
+ 5.201010000e-07 V_hig
+ 5.202000000e-07 V_hig
+ 5.202010000e-07 V_hig
+ 5.203000000e-07 V_hig
+ 5.203010000e-07 V_hig
+ 5.204000000e-07 V_hig
+ 5.204010000e-07 V_hig
+ 5.205000000e-07 V_hig
+ 5.205010000e-07 V_hig
+ 5.206000000e-07 V_hig
+ 5.206010000e-07 V_hig
+ 5.207000000e-07 V_hig
+ 5.207010000e-07 V_hig
+ 5.208000000e-07 V_hig
+ 5.208010000e-07 V_hig
+ 5.209000000e-07 V_hig
+ 5.209010000e-07 V_hig
+ 5.210000000e-07 V_hig
+ 5.210010000e-07 V_hig
+ 5.211000000e-07 V_hig
+ 5.211010000e-07 V_hig
+ 5.212000000e-07 V_hig
+ 5.212010000e-07 V_hig
+ 5.213000000e-07 V_hig
+ 5.213010000e-07 V_hig
+ 5.214000000e-07 V_hig
+ 5.214010000e-07 V_hig
+ 5.215000000e-07 V_hig
+ 5.215010000e-07 V_hig
+ 5.216000000e-07 V_hig
+ 5.216010000e-07 V_hig
+ 5.217000000e-07 V_hig
+ 5.217010000e-07 V_hig
+ 5.218000000e-07 V_hig
+ 5.218010000e-07 V_hig
+ 5.219000000e-07 V_hig
+ 5.219010000e-07 V_low
+ 5.220000000e-07 V_low
+ 5.220010000e-07 V_low
+ 5.221000000e-07 V_low
+ 5.221010000e-07 V_low
+ 5.222000000e-07 V_low
+ 5.222010000e-07 V_low
+ 5.223000000e-07 V_low
+ 5.223010000e-07 V_low
+ 5.224000000e-07 V_low
+ 5.224010000e-07 V_low
+ 5.225000000e-07 V_low
+ 5.225010000e-07 V_low
+ 5.226000000e-07 V_low
+ 5.226010000e-07 V_low
+ 5.227000000e-07 V_low
+ 5.227010000e-07 V_low
+ 5.228000000e-07 V_low
+ 5.228010000e-07 V_low
+ 5.229000000e-07 V_low
+ 5.229010000e-07 V_hig
+ 5.230000000e-07 V_hig
+ 5.230010000e-07 V_hig
+ 5.231000000e-07 V_hig
+ 5.231010000e-07 V_hig
+ 5.232000000e-07 V_hig
+ 5.232010000e-07 V_hig
+ 5.233000000e-07 V_hig
+ 5.233010000e-07 V_hig
+ 5.234000000e-07 V_hig
+ 5.234010000e-07 V_hig
+ 5.235000000e-07 V_hig
+ 5.235010000e-07 V_hig
+ 5.236000000e-07 V_hig
+ 5.236010000e-07 V_hig
+ 5.237000000e-07 V_hig
+ 5.237010000e-07 V_hig
+ 5.238000000e-07 V_hig
+ 5.238010000e-07 V_hig
+ 5.239000000e-07 V_hig
+ 5.239010000e-07 V_hig
+ 5.240000000e-07 V_hig
+ 5.240010000e-07 V_hig
+ 5.241000000e-07 V_hig
+ 5.241010000e-07 V_hig
+ 5.242000000e-07 V_hig
+ 5.242010000e-07 V_hig
+ 5.243000000e-07 V_hig
+ 5.243010000e-07 V_hig
+ 5.244000000e-07 V_hig
+ 5.244010000e-07 V_hig
+ 5.245000000e-07 V_hig
+ 5.245010000e-07 V_hig
+ 5.246000000e-07 V_hig
+ 5.246010000e-07 V_hig
+ 5.247000000e-07 V_hig
+ 5.247010000e-07 V_hig
+ 5.248000000e-07 V_hig
+ 5.248010000e-07 V_hig
+ 5.249000000e-07 V_hig
+ 5.249010000e-07 V_hig
+ 5.250000000e-07 V_hig
+ 5.250010000e-07 V_hig
+ 5.251000000e-07 V_hig
+ 5.251010000e-07 V_hig
+ 5.252000000e-07 V_hig
+ 5.252010000e-07 V_hig
+ 5.253000000e-07 V_hig
+ 5.253010000e-07 V_hig
+ 5.254000000e-07 V_hig
+ 5.254010000e-07 V_hig
+ 5.255000000e-07 V_hig
+ 5.255010000e-07 V_hig
+ 5.256000000e-07 V_hig
+ 5.256010000e-07 V_hig
+ 5.257000000e-07 V_hig
+ 5.257010000e-07 V_hig
+ 5.258000000e-07 V_hig
+ 5.258010000e-07 V_hig
+ 5.259000000e-07 V_hig
+ 5.259010000e-07 V_low
+ 5.260000000e-07 V_low
+ 5.260010000e-07 V_low
+ 5.261000000e-07 V_low
+ 5.261010000e-07 V_low
+ 5.262000000e-07 V_low
+ 5.262010000e-07 V_low
+ 5.263000000e-07 V_low
+ 5.263010000e-07 V_low
+ 5.264000000e-07 V_low
+ 5.264010000e-07 V_low
+ 5.265000000e-07 V_low
+ 5.265010000e-07 V_low
+ 5.266000000e-07 V_low
+ 5.266010000e-07 V_low
+ 5.267000000e-07 V_low
+ 5.267010000e-07 V_low
+ 5.268000000e-07 V_low
+ 5.268010000e-07 V_low
+ 5.269000000e-07 V_low
+ 5.269010000e-07 V_low
+ 5.270000000e-07 V_low
+ 5.270010000e-07 V_low
+ 5.271000000e-07 V_low
+ 5.271010000e-07 V_low
+ 5.272000000e-07 V_low
+ 5.272010000e-07 V_low
+ 5.273000000e-07 V_low
+ 5.273010000e-07 V_low
+ 5.274000000e-07 V_low
+ 5.274010000e-07 V_low
+ 5.275000000e-07 V_low
+ 5.275010000e-07 V_low
+ 5.276000000e-07 V_low
+ 5.276010000e-07 V_low
+ 5.277000000e-07 V_low
+ 5.277010000e-07 V_low
+ 5.278000000e-07 V_low
+ 5.278010000e-07 V_low
+ 5.279000000e-07 V_low
+ 5.279010000e-07 V_hig
+ 5.280000000e-07 V_hig
+ 5.280010000e-07 V_hig
+ 5.281000000e-07 V_hig
+ 5.281010000e-07 V_hig
+ 5.282000000e-07 V_hig
+ 5.282010000e-07 V_hig
+ 5.283000000e-07 V_hig
+ 5.283010000e-07 V_hig
+ 5.284000000e-07 V_hig
+ 5.284010000e-07 V_hig
+ 5.285000000e-07 V_hig
+ 5.285010000e-07 V_hig
+ 5.286000000e-07 V_hig
+ 5.286010000e-07 V_hig
+ 5.287000000e-07 V_hig
+ 5.287010000e-07 V_hig
+ 5.288000000e-07 V_hig
+ 5.288010000e-07 V_hig
+ 5.289000000e-07 V_hig
+ 5.289010000e-07 V_low
+ 5.290000000e-07 V_low
+ 5.290010000e-07 V_low
+ 5.291000000e-07 V_low
+ 5.291010000e-07 V_low
+ 5.292000000e-07 V_low
+ 5.292010000e-07 V_low
+ 5.293000000e-07 V_low
+ 5.293010000e-07 V_low
+ 5.294000000e-07 V_low
+ 5.294010000e-07 V_low
+ 5.295000000e-07 V_low
+ 5.295010000e-07 V_low
+ 5.296000000e-07 V_low
+ 5.296010000e-07 V_low
+ 5.297000000e-07 V_low
+ 5.297010000e-07 V_low
+ 5.298000000e-07 V_low
+ 5.298010000e-07 V_low
+ 5.299000000e-07 V_low
+ 5.299010000e-07 V_hig
+ 5.300000000e-07 V_hig
+ 5.300010000e-07 V_hig
+ 5.301000000e-07 V_hig
+ 5.301010000e-07 V_hig
+ 5.302000000e-07 V_hig
+ 5.302010000e-07 V_hig
+ 5.303000000e-07 V_hig
+ 5.303010000e-07 V_hig
+ 5.304000000e-07 V_hig
+ 5.304010000e-07 V_hig
+ 5.305000000e-07 V_hig
+ 5.305010000e-07 V_hig
+ 5.306000000e-07 V_hig
+ 5.306010000e-07 V_hig
+ 5.307000000e-07 V_hig
+ 5.307010000e-07 V_hig
+ 5.308000000e-07 V_hig
+ 5.308010000e-07 V_hig
+ 5.309000000e-07 V_hig
+ 5.309010000e-07 V_low
+ 5.310000000e-07 V_low
+ 5.310010000e-07 V_low
+ 5.311000000e-07 V_low
+ 5.311010000e-07 V_low
+ 5.312000000e-07 V_low
+ 5.312010000e-07 V_low
+ 5.313000000e-07 V_low
+ 5.313010000e-07 V_low
+ 5.314000000e-07 V_low
+ 5.314010000e-07 V_low
+ 5.315000000e-07 V_low
+ 5.315010000e-07 V_low
+ 5.316000000e-07 V_low
+ 5.316010000e-07 V_low
+ 5.317000000e-07 V_low
+ 5.317010000e-07 V_low
+ 5.318000000e-07 V_low
+ 5.318010000e-07 V_low
+ 5.319000000e-07 V_low
+ 5.319010000e-07 V_low
+ 5.320000000e-07 V_low
+ 5.320010000e-07 V_low
+ 5.321000000e-07 V_low
+ 5.321010000e-07 V_low
+ 5.322000000e-07 V_low
+ 5.322010000e-07 V_low
+ 5.323000000e-07 V_low
+ 5.323010000e-07 V_low
+ 5.324000000e-07 V_low
+ 5.324010000e-07 V_low
+ 5.325000000e-07 V_low
+ 5.325010000e-07 V_low
+ 5.326000000e-07 V_low
+ 5.326010000e-07 V_low
+ 5.327000000e-07 V_low
+ 5.327010000e-07 V_low
+ 5.328000000e-07 V_low
+ 5.328010000e-07 V_low
+ 5.329000000e-07 V_low
+ 5.329010000e-07 V_low
+ 5.330000000e-07 V_low
+ 5.330010000e-07 V_low
+ 5.331000000e-07 V_low
+ 5.331010000e-07 V_low
+ 5.332000000e-07 V_low
+ 5.332010000e-07 V_low
+ 5.333000000e-07 V_low
+ 5.333010000e-07 V_low
+ 5.334000000e-07 V_low
+ 5.334010000e-07 V_low
+ 5.335000000e-07 V_low
+ 5.335010000e-07 V_low
+ 5.336000000e-07 V_low
+ 5.336010000e-07 V_low
+ 5.337000000e-07 V_low
+ 5.337010000e-07 V_low
+ 5.338000000e-07 V_low
+ 5.338010000e-07 V_low
+ 5.339000000e-07 V_low
+ 5.339010000e-07 V_hig
+ 5.340000000e-07 V_hig
+ 5.340010000e-07 V_hig
+ 5.341000000e-07 V_hig
+ 5.341010000e-07 V_hig
+ 5.342000000e-07 V_hig
+ 5.342010000e-07 V_hig
+ 5.343000000e-07 V_hig
+ 5.343010000e-07 V_hig
+ 5.344000000e-07 V_hig
+ 5.344010000e-07 V_hig
+ 5.345000000e-07 V_hig
+ 5.345010000e-07 V_hig
+ 5.346000000e-07 V_hig
+ 5.346010000e-07 V_hig
+ 5.347000000e-07 V_hig
+ 5.347010000e-07 V_hig
+ 5.348000000e-07 V_hig
+ 5.348010000e-07 V_hig
+ 5.349000000e-07 V_hig
+ 5.349010000e-07 V_low
+ 5.350000000e-07 V_low
+ 5.350010000e-07 V_low
+ 5.351000000e-07 V_low
+ 5.351010000e-07 V_low
+ 5.352000000e-07 V_low
+ 5.352010000e-07 V_low
+ 5.353000000e-07 V_low
+ 5.353010000e-07 V_low
+ 5.354000000e-07 V_low
+ 5.354010000e-07 V_low
+ 5.355000000e-07 V_low
+ 5.355010000e-07 V_low
+ 5.356000000e-07 V_low
+ 5.356010000e-07 V_low
+ 5.357000000e-07 V_low
+ 5.357010000e-07 V_low
+ 5.358000000e-07 V_low
+ 5.358010000e-07 V_low
+ 5.359000000e-07 V_low
+ 5.359010000e-07 V_low
+ 5.360000000e-07 V_low
+ 5.360010000e-07 V_low
+ 5.361000000e-07 V_low
+ 5.361010000e-07 V_low
+ 5.362000000e-07 V_low
+ 5.362010000e-07 V_low
+ 5.363000000e-07 V_low
+ 5.363010000e-07 V_low
+ 5.364000000e-07 V_low
+ 5.364010000e-07 V_low
+ 5.365000000e-07 V_low
+ 5.365010000e-07 V_low
+ 5.366000000e-07 V_low
+ 5.366010000e-07 V_low
+ 5.367000000e-07 V_low
+ 5.367010000e-07 V_low
+ 5.368000000e-07 V_low
+ 5.368010000e-07 V_low
+ 5.369000000e-07 V_low
+ 5.369010000e-07 V_hig
+ 5.370000000e-07 V_hig
+ 5.370010000e-07 V_hig
+ 5.371000000e-07 V_hig
+ 5.371010000e-07 V_hig
+ 5.372000000e-07 V_hig
+ 5.372010000e-07 V_hig
+ 5.373000000e-07 V_hig
+ 5.373010000e-07 V_hig
+ 5.374000000e-07 V_hig
+ 5.374010000e-07 V_hig
+ 5.375000000e-07 V_hig
+ 5.375010000e-07 V_hig
+ 5.376000000e-07 V_hig
+ 5.376010000e-07 V_hig
+ 5.377000000e-07 V_hig
+ 5.377010000e-07 V_hig
+ 5.378000000e-07 V_hig
+ 5.378010000e-07 V_hig
+ 5.379000000e-07 V_hig
+ 5.379010000e-07 V_low
+ 5.380000000e-07 V_low
+ 5.380010000e-07 V_low
+ 5.381000000e-07 V_low
+ 5.381010000e-07 V_low
+ 5.382000000e-07 V_low
+ 5.382010000e-07 V_low
+ 5.383000000e-07 V_low
+ 5.383010000e-07 V_low
+ 5.384000000e-07 V_low
+ 5.384010000e-07 V_low
+ 5.385000000e-07 V_low
+ 5.385010000e-07 V_low
+ 5.386000000e-07 V_low
+ 5.386010000e-07 V_low
+ 5.387000000e-07 V_low
+ 5.387010000e-07 V_low
+ 5.388000000e-07 V_low
+ 5.388010000e-07 V_low
+ 5.389000000e-07 V_low
+ 5.389010000e-07 V_low
+ 5.390000000e-07 V_low
+ 5.390010000e-07 V_low
+ 5.391000000e-07 V_low
+ 5.391010000e-07 V_low
+ 5.392000000e-07 V_low
+ 5.392010000e-07 V_low
+ 5.393000000e-07 V_low
+ 5.393010000e-07 V_low
+ 5.394000000e-07 V_low
+ 5.394010000e-07 V_low
+ 5.395000000e-07 V_low
+ 5.395010000e-07 V_low
+ 5.396000000e-07 V_low
+ 5.396010000e-07 V_low
+ 5.397000000e-07 V_low
+ 5.397010000e-07 V_low
+ 5.398000000e-07 V_low
+ 5.398010000e-07 V_low
+ 5.399000000e-07 V_low
+ 5.399010000e-07 V_low
+ 5.400000000e-07 V_low
+ 5.400010000e-07 V_low
+ 5.401000000e-07 V_low
+ 5.401010000e-07 V_low
+ 5.402000000e-07 V_low
+ 5.402010000e-07 V_low
+ 5.403000000e-07 V_low
+ 5.403010000e-07 V_low
+ 5.404000000e-07 V_low
+ 5.404010000e-07 V_low
+ 5.405000000e-07 V_low
+ 5.405010000e-07 V_low
+ 5.406000000e-07 V_low
+ 5.406010000e-07 V_low
+ 5.407000000e-07 V_low
+ 5.407010000e-07 V_low
+ 5.408000000e-07 V_low
+ 5.408010000e-07 V_low
+ 5.409000000e-07 V_low
+ 5.409010000e-07 V_hig
+ 5.410000000e-07 V_hig
+ 5.410010000e-07 V_hig
+ 5.411000000e-07 V_hig
+ 5.411010000e-07 V_hig
+ 5.412000000e-07 V_hig
+ 5.412010000e-07 V_hig
+ 5.413000000e-07 V_hig
+ 5.413010000e-07 V_hig
+ 5.414000000e-07 V_hig
+ 5.414010000e-07 V_hig
+ 5.415000000e-07 V_hig
+ 5.415010000e-07 V_hig
+ 5.416000000e-07 V_hig
+ 5.416010000e-07 V_hig
+ 5.417000000e-07 V_hig
+ 5.417010000e-07 V_hig
+ 5.418000000e-07 V_hig
+ 5.418010000e-07 V_hig
+ 5.419000000e-07 V_hig
+ 5.419010000e-07 V_low
+ 5.420000000e-07 V_low
+ 5.420010000e-07 V_low
+ 5.421000000e-07 V_low
+ 5.421010000e-07 V_low
+ 5.422000000e-07 V_low
+ 5.422010000e-07 V_low
+ 5.423000000e-07 V_low
+ 5.423010000e-07 V_low
+ 5.424000000e-07 V_low
+ 5.424010000e-07 V_low
+ 5.425000000e-07 V_low
+ 5.425010000e-07 V_low
+ 5.426000000e-07 V_low
+ 5.426010000e-07 V_low
+ 5.427000000e-07 V_low
+ 5.427010000e-07 V_low
+ 5.428000000e-07 V_low
+ 5.428010000e-07 V_low
+ 5.429000000e-07 V_low
+ 5.429010000e-07 V_low
+ 5.430000000e-07 V_low
+ 5.430010000e-07 V_low
+ 5.431000000e-07 V_low
+ 5.431010000e-07 V_low
+ 5.432000000e-07 V_low
+ 5.432010000e-07 V_low
+ 5.433000000e-07 V_low
+ 5.433010000e-07 V_low
+ 5.434000000e-07 V_low
+ 5.434010000e-07 V_low
+ 5.435000000e-07 V_low
+ 5.435010000e-07 V_low
+ 5.436000000e-07 V_low
+ 5.436010000e-07 V_low
+ 5.437000000e-07 V_low
+ 5.437010000e-07 V_low
+ 5.438000000e-07 V_low
+ 5.438010000e-07 V_low
+ 5.439000000e-07 V_low
+ 5.439010000e-07 V_low
+ 5.440000000e-07 V_low
+ 5.440010000e-07 V_low
+ 5.441000000e-07 V_low
+ 5.441010000e-07 V_low
+ 5.442000000e-07 V_low
+ 5.442010000e-07 V_low
+ 5.443000000e-07 V_low
+ 5.443010000e-07 V_low
+ 5.444000000e-07 V_low
+ 5.444010000e-07 V_low
+ 5.445000000e-07 V_low
+ 5.445010000e-07 V_low
+ 5.446000000e-07 V_low
+ 5.446010000e-07 V_low
+ 5.447000000e-07 V_low
+ 5.447010000e-07 V_low
+ 5.448000000e-07 V_low
+ 5.448010000e-07 V_low
+ 5.449000000e-07 V_low
+ 5.449010000e-07 V_hig
+ 5.450000000e-07 V_hig
+ 5.450010000e-07 V_hig
+ 5.451000000e-07 V_hig
+ 5.451010000e-07 V_hig
+ 5.452000000e-07 V_hig
+ 5.452010000e-07 V_hig
+ 5.453000000e-07 V_hig
+ 5.453010000e-07 V_hig
+ 5.454000000e-07 V_hig
+ 5.454010000e-07 V_hig
+ 5.455000000e-07 V_hig
+ 5.455010000e-07 V_hig
+ 5.456000000e-07 V_hig
+ 5.456010000e-07 V_hig
+ 5.457000000e-07 V_hig
+ 5.457010000e-07 V_hig
+ 5.458000000e-07 V_hig
+ 5.458010000e-07 V_hig
+ 5.459000000e-07 V_hig
+ 5.459010000e-07 V_low
+ 5.460000000e-07 V_low
+ 5.460010000e-07 V_low
+ 5.461000000e-07 V_low
+ 5.461010000e-07 V_low
+ 5.462000000e-07 V_low
+ 5.462010000e-07 V_low
+ 5.463000000e-07 V_low
+ 5.463010000e-07 V_low
+ 5.464000000e-07 V_low
+ 5.464010000e-07 V_low
+ 5.465000000e-07 V_low
+ 5.465010000e-07 V_low
+ 5.466000000e-07 V_low
+ 5.466010000e-07 V_low
+ 5.467000000e-07 V_low
+ 5.467010000e-07 V_low
+ 5.468000000e-07 V_low
+ 5.468010000e-07 V_low
+ 5.469000000e-07 V_low
+ 5.469010000e-07 V_hig
+ 5.470000000e-07 V_hig
+ 5.470010000e-07 V_hig
+ 5.471000000e-07 V_hig
+ 5.471010000e-07 V_hig
+ 5.472000000e-07 V_hig
+ 5.472010000e-07 V_hig
+ 5.473000000e-07 V_hig
+ 5.473010000e-07 V_hig
+ 5.474000000e-07 V_hig
+ 5.474010000e-07 V_hig
+ 5.475000000e-07 V_hig
+ 5.475010000e-07 V_hig
+ 5.476000000e-07 V_hig
+ 5.476010000e-07 V_hig
+ 5.477000000e-07 V_hig
+ 5.477010000e-07 V_hig
+ 5.478000000e-07 V_hig
+ 5.478010000e-07 V_hig
+ 5.479000000e-07 V_hig
+ 5.479010000e-07 V_low
+ 5.480000000e-07 V_low
+ 5.480010000e-07 V_low
+ 5.481000000e-07 V_low
+ 5.481010000e-07 V_low
+ 5.482000000e-07 V_low
+ 5.482010000e-07 V_low
+ 5.483000000e-07 V_low
+ 5.483010000e-07 V_low
+ 5.484000000e-07 V_low
+ 5.484010000e-07 V_low
+ 5.485000000e-07 V_low
+ 5.485010000e-07 V_low
+ 5.486000000e-07 V_low
+ 5.486010000e-07 V_low
+ 5.487000000e-07 V_low
+ 5.487010000e-07 V_low
+ 5.488000000e-07 V_low
+ 5.488010000e-07 V_low
+ 5.489000000e-07 V_low
+ 5.489010000e-07 V_low
+ 5.490000000e-07 V_low
+ 5.490010000e-07 V_low
+ 5.491000000e-07 V_low
+ 5.491010000e-07 V_low
+ 5.492000000e-07 V_low
+ 5.492010000e-07 V_low
+ 5.493000000e-07 V_low
+ 5.493010000e-07 V_low
+ 5.494000000e-07 V_low
+ 5.494010000e-07 V_low
+ 5.495000000e-07 V_low
+ 5.495010000e-07 V_low
+ 5.496000000e-07 V_low
+ 5.496010000e-07 V_low
+ 5.497000000e-07 V_low
+ 5.497010000e-07 V_low
+ 5.498000000e-07 V_low
+ 5.498010000e-07 V_low
+ 5.499000000e-07 V_low
+ 5.499010000e-07 V_hig
+ 5.500000000e-07 V_hig
+ 5.500010000e-07 V_hig
+ 5.501000000e-07 V_hig
+ 5.501010000e-07 V_hig
+ 5.502000000e-07 V_hig
+ 5.502010000e-07 V_hig
+ 5.503000000e-07 V_hig
+ 5.503010000e-07 V_hig
+ 5.504000000e-07 V_hig
+ 5.504010000e-07 V_hig
+ 5.505000000e-07 V_hig
+ 5.505010000e-07 V_hig
+ 5.506000000e-07 V_hig
+ 5.506010000e-07 V_hig
+ 5.507000000e-07 V_hig
+ 5.507010000e-07 V_hig
+ 5.508000000e-07 V_hig
+ 5.508010000e-07 V_hig
+ 5.509000000e-07 V_hig
+ 5.509010000e-07 V_hig
+ 5.510000000e-07 V_hig
+ 5.510010000e-07 V_hig
+ 5.511000000e-07 V_hig
+ 5.511010000e-07 V_hig
+ 5.512000000e-07 V_hig
+ 5.512010000e-07 V_hig
+ 5.513000000e-07 V_hig
+ 5.513010000e-07 V_hig
+ 5.514000000e-07 V_hig
+ 5.514010000e-07 V_hig
+ 5.515000000e-07 V_hig
+ 5.515010000e-07 V_hig
+ 5.516000000e-07 V_hig
+ 5.516010000e-07 V_hig
+ 5.517000000e-07 V_hig
+ 5.517010000e-07 V_hig
+ 5.518000000e-07 V_hig
+ 5.518010000e-07 V_hig
+ 5.519000000e-07 V_hig
+ 5.519010000e-07 V_low
+ 5.520000000e-07 V_low
+ 5.520010000e-07 V_low
+ 5.521000000e-07 V_low
+ 5.521010000e-07 V_low
+ 5.522000000e-07 V_low
+ 5.522010000e-07 V_low
+ 5.523000000e-07 V_low
+ 5.523010000e-07 V_low
+ 5.524000000e-07 V_low
+ 5.524010000e-07 V_low
+ 5.525000000e-07 V_low
+ 5.525010000e-07 V_low
+ 5.526000000e-07 V_low
+ 5.526010000e-07 V_low
+ 5.527000000e-07 V_low
+ 5.527010000e-07 V_low
+ 5.528000000e-07 V_low
+ 5.528010000e-07 V_low
+ 5.529000000e-07 V_low
+ 5.529010000e-07 V_low
+ 5.530000000e-07 V_low
+ 5.530010000e-07 V_low
+ 5.531000000e-07 V_low
+ 5.531010000e-07 V_low
+ 5.532000000e-07 V_low
+ 5.532010000e-07 V_low
+ 5.533000000e-07 V_low
+ 5.533010000e-07 V_low
+ 5.534000000e-07 V_low
+ 5.534010000e-07 V_low
+ 5.535000000e-07 V_low
+ 5.535010000e-07 V_low
+ 5.536000000e-07 V_low
+ 5.536010000e-07 V_low
+ 5.537000000e-07 V_low
+ 5.537010000e-07 V_low
+ 5.538000000e-07 V_low
+ 5.538010000e-07 V_low
+ 5.539000000e-07 V_low
+ 5.539010000e-07 V_low
+ 5.540000000e-07 V_low
+ 5.540010000e-07 V_low
+ 5.541000000e-07 V_low
+ 5.541010000e-07 V_low
+ 5.542000000e-07 V_low
+ 5.542010000e-07 V_low
+ 5.543000000e-07 V_low
+ 5.543010000e-07 V_low
+ 5.544000000e-07 V_low
+ 5.544010000e-07 V_low
+ 5.545000000e-07 V_low
+ 5.545010000e-07 V_low
+ 5.546000000e-07 V_low
+ 5.546010000e-07 V_low
+ 5.547000000e-07 V_low
+ 5.547010000e-07 V_low
+ 5.548000000e-07 V_low
+ 5.548010000e-07 V_low
+ 5.549000000e-07 V_low
+ 5.549010000e-07 V_low
+ 5.550000000e-07 V_low
+ 5.550010000e-07 V_low
+ 5.551000000e-07 V_low
+ 5.551010000e-07 V_low
+ 5.552000000e-07 V_low
+ 5.552010000e-07 V_low
+ 5.553000000e-07 V_low
+ 5.553010000e-07 V_low
+ 5.554000000e-07 V_low
+ 5.554010000e-07 V_low
+ 5.555000000e-07 V_low
+ 5.555010000e-07 V_low
+ 5.556000000e-07 V_low
+ 5.556010000e-07 V_low
+ 5.557000000e-07 V_low
+ 5.557010000e-07 V_low
+ 5.558000000e-07 V_low
+ 5.558010000e-07 V_low
+ 5.559000000e-07 V_low
+ 5.559010000e-07 V_low
+ 5.560000000e-07 V_low
+ 5.560010000e-07 V_low
+ 5.561000000e-07 V_low
+ 5.561010000e-07 V_low
+ 5.562000000e-07 V_low
+ 5.562010000e-07 V_low
+ 5.563000000e-07 V_low
+ 5.563010000e-07 V_low
+ 5.564000000e-07 V_low
+ 5.564010000e-07 V_low
+ 5.565000000e-07 V_low
+ 5.565010000e-07 V_low
+ 5.566000000e-07 V_low
+ 5.566010000e-07 V_low
+ 5.567000000e-07 V_low
+ 5.567010000e-07 V_low
+ 5.568000000e-07 V_low
+ 5.568010000e-07 V_low
+ 5.569000000e-07 V_low
+ 5.569010000e-07 V_low
+ 5.570000000e-07 V_low
+ 5.570010000e-07 V_low
+ 5.571000000e-07 V_low
+ 5.571010000e-07 V_low
+ 5.572000000e-07 V_low
+ 5.572010000e-07 V_low
+ 5.573000000e-07 V_low
+ 5.573010000e-07 V_low
+ 5.574000000e-07 V_low
+ 5.574010000e-07 V_low
+ 5.575000000e-07 V_low
+ 5.575010000e-07 V_low
+ 5.576000000e-07 V_low
+ 5.576010000e-07 V_low
+ 5.577000000e-07 V_low
+ 5.577010000e-07 V_low
+ 5.578000000e-07 V_low
+ 5.578010000e-07 V_low
+ 5.579000000e-07 V_low
+ 5.579010000e-07 V_hig
+ 5.580000000e-07 V_hig
+ 5.580010000e-07 V_hig
+ 5.581000000e-07 V_hig
+ 5.581010000e-07 V_hig
+ 5.582000000e-07 V_hig
+ 5.582010000e-07 V_hig
+ 5.583000000e-07 V_hig
+ 5.583010000e-07 V_hig
+ 5.584000000e-07 V_hig
+ 5.584010000e-07 V_hig
+ 5.585000000e-07 V_hig
+ 5.585010000e-07 V_hig
+ 5.586000000e-07 V_hig
+ 5.586010000e-07 V_hig
+ 5.587000000e-07 V_hig
+ 5.587010000e-07 V_hig
+ 5.588000000e-07 V_hig
+ 5.588010000e-07 V_hig
+ 5.589000000e-07 V_hig
+ 5.589010000e-07 V_hig
+ 5.590000000e-07 V_hig
+ 5.590010000e-07 V_hig
+ 5.591000000e-07 V_hig
+ 5.591010000e-07 V_hig
+ 5.592000000e-07 V_hig
+ 5.592010000e-07 V_hig
+ 5.593000000e-07 V_hig
+ 5.593010000e-07 V_hig
+ 5.594000000e-07 V_hig
+ 5.594010000e-07 V_hig
+ 5.595000000e-07 V_hig
+ 5.595010000e-07 V_hig
+ 5.596000000e-07 V_hig
+ 5.596010000e-07 V_hig
+ 5.597000000e-07 V_hig
+ 5.597010000e-07 V_hig
+ 5.598000000e-07 V_hig
+ 5.598010000e-07 V_hig
+ 5.599000000e-07 V_hig
+ 5.599010000e-07 V_hig
+ 5.600000000e-07 V_hig
+ 5.600010000e-07 V_hig
+ 5.601000000e-07 V_hig
+ 5.601010000e-07 V_hig
+ 5.602000000e-07 V_hig
+ 5.602010000e-07 V_hig
+ 5.603000000e-07 V_hig
+ 5.603010000e-07 V_hig
+ 5.604000000e-07 V_hig
+ 5.604010000e-07 V_hig
+ 5.605000000e-07 V_hig
+ 5.605010000e-07 V_hig
+ 5.606000000e-07 V_hig
+ 5.606010000e-07 V_hig
+ 5.607000000e-07 V_hig
+ 5.607010000e-07 V_hig
+ 5.608000000e-07 V_hig
+ 5.608010000e-07 V_hig
+ 5.609000000e-07 V_hig
+ 5.609010000e-07 V_low
+ 5.610000000e-07 V_low
+ 5.610010000e-07 V_low
+ 5.611000000e-07 V_low
+ 5.611010000e-07 V_low
+ 5.612000000e-07 V_low
+ 5.612010000e-07 V_low
+ 5.613000000e-07 V_low
+ 5.613010000e-07 V_low
+ 5.614000000e-07 V_low
+ 5.614010000e-07 V_low
+ 5.615000000e-07 V_low
+ 5.615010000e-07 V_low
+ 5.616000000e-07 V_low
+ 5.616010000e-07 V_low
+ 5.617000000e-07 V_low
+ 5.617010000e-07 V_low
+ 5.618000000e-07 V_low
+ 5.618010000e-07 V_low
+ 5.619000000e-07 V_low
+ 5.619010000e-07 V_low
+ 5.620000000e-07 V_low
+ 5.620010000e-07 V_low
+ 5.621000000e-07 V_low
+ 5.621010000e-07 V_low
+ 5.622000000e-07 V_low
+ 5.622010000e-07 V_low
+ 5.623000000e-07 V_low
+ 5.623010000e-07 V_low
+ 5.624000000e-07 V_low
+ 5.624010000e-07 V_low
+ 5.625000000e-07 V_low
+ 5.625010000e-07 V_low
+ 5.626000000e-07 V_low
+ 5.626010000e-07 V_low
+ 5.627000000e-07 V_low
+ 5.627010000e-07 V_low
+ 5.628000000e-07 V_low
+ 5.628010000e-07 V_low
+ 5.629000000e-07 V_low
+ 5.629010000e-07 V_hig
+ 5.630000000e-07 V_hig
+ 5.630010000e-07 V_hig
+ 5.631000000e-07 V_hig
+ 5.631010000e-07 V_hig
+ 5.632000000e-07 V_hig
+ 5.632010000e-07 V_hig
+ 5.633000000e-07 V_hig
+ 5.633010000e-07 V_hig
+ 5.634000000e-07 V_hig
+ 5.634010000e-07 V_hig
+ 5.635000000e-07 V_hig
+ 5.635010000e-07 V_hig
+ 5.636000000e-07 V_hig
+ 5.636010000e-07 V_hig
+ 5.637000000e-07 V_hig
+ 5.637010000e-07 V_hig
+ 5.638000000e-07 V_hig
+ 5.638010000e-07 V_hig
+ 5.639000000e-07 V_hig
+ 5.639010000e-07 V_low
+ 5.640000000e-07 V_low
+ 5.640010000e-07 V_low
+ 5.641000000e-07 V_low
+ 5.641010000e-07 V_low
+ 5.642000000e-07 V_low
+ 5.642010000e-07 V_low
+ 5.643000000e-07 V_low
+ 5.643010000e-07 V_low
+ 5.644000000e-07 V_low
+ 5.644010000e-07 V_low
+ 5.645000000e-07 V_low
+ 5.645010000e-07 V_low
+ 5.646000000e-07 V_low
+ 5.646010000e-07 V_low
+ 5.647000000e-07 V_low
+ 5.647010000e-07 V_low
+ 5.648000000e-07 V_low
+ 5.648010000e-07 V_low
+ 5.649000000e-07 V_low
+ 5.649010000e-07 V_low
+ 5.650000000e-07 V_low
+ 5.650010000e-07 V_low
+ 5.651000000e-07 V_low
+ 5.651010000e-07 V_low
+ 5.652000000e-07 V_low
+ 5.652010000e-07 V_low
+ 5.653000000e-07 V_low
+ 5.653010000e-07 V_low
+ 5.654000000e-07 V_low
+ 5.654010000e-07 V_low
+ 5.655000000e-07 V_low
+ 5.655010000e-07 V_low
+ 5.656000000e-07 V_low
+ 5.656010000e-07 V_low
+ 5.657000000e-07 V_low
+ 5.657010000e-07 V_low
+ 5.658000000e-07 V_low
+ 5.658010000e-07 V_low
+ 5.659000000e-07 V_low
+ 5.659010000e-07 V_hig
+ 5.660000000e-07 V_hig
+ 5.660010000e-07 V_hig
+ 5.661000000e-07 V_hig
+ 5.661010000e-07 V_hig
+ 5.662000000e-07 V_hig
+ 5.662010000e-07 V_hig
+ 5.663000000e-07 V_hig
+ 5.663010000e-07 V_hig
+ 5.664000000e-07 V_hig
+ 5.664010000e-07 V_hig
+ 5.665000000e-07 V_hig
+ 5.665010000e-07 V_hig
+ 5.666000000e-07 V_hig
+ 5.666010000e-07 V_hig
+ 5.667000000e-07 V_hig
+ 5.667010000e-07 V_hig
+ 5.668000000e-07 V_hig
+ 5.668010000e-07 V_hig
+ 5.669000000e-07 V_hig
+ 5.669010000e-07 V_low
+ 5.670000000e-07 V_low
+ 5.670010000e-07 V_low
+ 5.671000000e-07 V_low
+ 5.671010000e-07 V_low
+ 5.672000000e-07 V_low
+ 5.672010000e-07 V_low
+ 5.673000000e-07 V_low
+ 5.673010000e-07 V_low
+ 5.674000000e-07 V_low
+ 5.674010000e-07 V_low
+ 5.675000000e-07 V_low
+ 5.675010000e-07 V_low
+ 5.676000000e-07 V_low
+ 5.676010000e-07 V_low
+ 5.677000000e-07 V_low
+ 5.677010000e-07 V_low
+ 5.678000000e-07 V_low
+ 5.678010000e-07 V_low
+ 5.679000000e-07 V_low
+ 5.679010000e-07 V_low
+ 5.680000000e-07 V_low
+ 5.680010000e-07 V_low
+ 5.681000000e-07 V_low
+ 5.681010000e-07 V_low
+ 5.682000000e-07 V_low
+ 5.682010000e-07 V_low
+ 5.683000000e-07 V_low
+ 5.683010000e-07 V_low
+ 5.684000000e-07 V_low
+ 5.684010000e-07 V_low
+ 5.685000000e-07 V_low
+ 5.685010000e-07 V_low
+ 5.686000000e-07 V_low
+ 5.686010000e-07 V_low
+ 5.687000000e-07 V_low
+ 5.687010000e-07 V_low
+ 5.688000000e-07 V_low
+ 5.688010000e-07 V_low
+ 5.689000000e-07 V_low
+ 5.689010000e-07 V_low
+ 5.690000000e-07 V_low
+ 5.690010000e-07 V_low
+ 5.691000000e-07 V_low
+ 5.691010000e-07 V_low
+ 5.692000000e-07 V_low
+ 5.692010000e-07 V_low
+ 5.693000000e-07 V_low
+ 5.693010000e-07 V_low
+ 5.694000000e-07 V_low
+ 5.694010000e-07 V_low
+ 5.695000000e-07 V_low
+ 5.695010000e-07 V_low
+ 5.696000000e-07 V_low
+ 5.696010000e-07 V_low
+ 5.697000000e-07 V_low
+ 5.697010000e-07 V_low
+ 5.698000000e-07 V_low
+ 5.698010000e-07 V_low
+ 5.699000000e-07 V_low
+ 5.699010000e-07 V_low
+ 5.700000000e-07 V_low
+ 5.700010000e-07 V_low
+ 5.701000000e-07 V_low
+ 5.701010000e-07 V_low
+ 5.702000000e-07 V_low
+ 5.702010000e-07 V_low
+ 5.703000000e-07 V_low
+ 5.703010000e-07 V_low
+ 5.704000000e-07 V_low
+ 5.704010000e-07 V_low
+ 5.705000000e-07 V_low
+ 5.705010000e-07 V_low
+ 5.706000000e-07 V_low
+ 5.706010000e-07 V_low
+ 5.707000000e-07 V_low
+ 5.707010000e-07 V_low
+ 5.708000000e-07 V_low
+ 5.708010000e-07 V_low
+ 5.709000000e-07 V_low
+ 5.709010000e-07 V_low
+ 5.710000000e-07 V_low
+ 5.710010000e-07 V_low
+ 5.711000000e-07 V_low
+ 5.711010000e-07 V_low
+ 5.712000000e-07 V_low
+ 5.712010000e-07 V_low
+ 5.713000000e-07 V_low
+ 5.713010000e-07 V_low
+ 5.714000000e-07 V_low
+ 5.714010000e-07 V_low
+ 5.715000000e-07 V_low
+ 5.715010000e-07 V_low
+ 5.716000000e-07 V_low
+ 5.716010000e-07 V_low
+ 5.717000000e-07 V_low
+ 5.717010000e-07 V_low
+ 5.718000000e-07 V_low
+ 5.718010000e-07 V_low
+ 5.719000000e-07 V_low
+ 5.719010000e-07 V_hig
+ 5.720000000e-07 V_hig
+ 5.720010000e-07 V_hig
+ 5.721000000e-07 V_hig
+ 5.721010000e-07 V_hig
+ 5.722000000e-07 V_hig
+ 5.722010000e-07 V_hig
+ 5.723000000e-07 V_hig
+ 5.723010000e-07 V_hig
+ 5.724000000e-07 V_hig
+ 5.724010000e-07 V_hig
+ 5.725000000e-07 V_hig
+ 5.725010000e-07 V_hig
+ 5.726000000e-07 V_hig
+ 5.726010000e-07 V_hig
+ 5.727000000e-07 V_hig
+ 5.727010000e-07 V_hig
+ 5.728000000e-07 V_hig
+ 5.728010000e-07 V_hig
+ 5.729000000e-07 V_hig
+ 5.729010000e-07 V_low
+ 5.730000000e-07 V_low
+ 5.730010000e-07 V_low
+ 5.731000000e-07 V_low
+ 5.731010000e-07 V_low
+ 5.732000000e-07 V_low
+ 5.732010000e-07 V_low
+ 5.733000000e-07 V_low
+ 5.733010000e-07 V_low
+ 5.734000000e-07 V_low
+ 5.734010000e-07 V_low
+ 5.735000000e-07 V_low
+ 5.735010000e-07 V_low
+ 5.736000000e-07 V_low
+ 5.736010000e-07 V_low
+ 5.737000000e-07 V_low
+ 5.737010000e-07 V_low
+ 5.738000000e-07 V_low
+ 5.738010000e-07 V_low
+ 5.739000000e-07 V_low
+ 5.739010000e-07 V_hig
+ 5.740000000e-07 V_hig
+ 5.740010000e-07 V_hig
+ 5.741000000e-07 V_hig
+ 5.741010000e-07 V_hig
+ 5.742000000e-07 V_hig
+ 5.742010000e-07 V_hig
+ 5.743000000e-07 V_hig
+ 5.743010000e-07 V_hig
+ 5.744000000e-07 V_hig
+ 5.744010000e-07 V_hig
+ 5.745000000e-07 V_hig
+ 5.745010000e-07 V_hig
+ 5.746000000e-07 V_hig
+ 5.746010000e-07 V_hig
+ 5.747000000e-07 V_hig
+ 5.747010000e-07 V_hig
+ 5.748000000e-07 V_hig
+ 5.748010000e-07 V_hig
+ 5.749000000e-07 V_hig
+ 5.749010000e-07 V_low
+ 5.750000000e-07 V_low
+ 5.750010000e-07 V_low
+ 5.751000000e-07 V_low
+ 5.751010000e-07 V_low
+ 5.752000000e-07 V_low
+ 5.752010000e-07 V_low
+ 5.753000000e-07 V_low
+ 5.753010000e-07 V_low
+ 5.754000000e-07 V_low
+ 5.754010000e-07 V_low
+ 5.755000000e-07 V_low
+ 5.755010000e-07 V_low
+ 5.756000000e-07 V_low
+ 5.756010000e-07 V_low
+ 5.757000000e-07 V_low
+ 5.757010000e-07 V_low
+ 5.758000000e-07 V_low
+ 5.758010000e-07 V_low
+ 5.759000000e-07 V_low
+ 5.759010000e-07 V_hig
+ 5.760000000e-07 V_hig
+ 5.760010000e-07 V_hig
+ 5.761000000e-07 V_hig
+ 5.761010000e-07 V_hig
+ 5.762000000e-07 V_hig
+ 5.762010000e-07 V_hig
+ 5.763000000e-07 V_hig
+ 5.763010000e-07 V_hig
+ 5.764000000e-07 V_hig
+ 5.764010000e-07 V_hig
+ 5.765000000e-07 V_hig
+ 5.765010000e-07 V_hig
+ 5.766000000e-07 V_hig
+ 5.766010000e-07 V_hig
+ 5.767000000e-07 V_hig
+ 5.767010000e-07 V_hig
+ 5.768000000e-07 V_hig
+ 5.768010000e-07 V_hig
+ 5.769000000e-07 V_hig
+ 5.769010000e-07 V_low
+ 5.770000000e-07 V_low
+ 5.770010000e-07 V_low
+ 5.771000000e-07 V_low
+ 5.771010000e-07 V_low
+ 5.772000000e-07 V_low
+ 5.772010000e-07 V_low
+ 5.773000000e-07 V_low
+ 5.773010000e-07 V_low
+ 5.774000000e-07 V_low
+ 5.774010000e-07 V_low
+ 5.775000000e-07 V_low
+ 5.775010000e-07 V_low
+ 5.776000000e-07 V_low
+ 5.776010000e-07 V_low
+ 5.777000000e-07 V_low
+ 5.777010000e-07 V_low
+ 5.778000000e-07 V_low
+ 5.778010000e-07 V_low
+ 5.779000000e-07 V_low
+ 5.779010000e-07 V_low
+ 5.780000000e-07 V_low
+ 5.780010000e-07 V_low
+ 5.781000000e-07 V_low
+ 5.781010000e-07 V_low
+ 5.782000000e-07 V_low
+ 5.782010000e-07 V_low
+ 5.783000000e-07 V_low
+ 5.783010000e-07 V_low
+ 5.784000000e-07 V_low
+ 5.784010000e-07 V_low
+ 5.785000000e-07 V_low
+ 5.785010000e-07 V_low
+ 5.786000000e-07 V_low
+ 5.786010000e-07 V_low
+ 5.787000000e-07 V_low
+ 5.787010000e-07 V_low
+ 5.788000000e-07 V_low
+ 5.788010000e-07 V_low
+ 5.789000000e-07 V_low
+ 5.789010000e-07 V_hig
+ 5.790000000e-07 V_hig
+ 5.790010000e-07 V_hig
+ 5.791000000e-07 V_hig
+ 5.791010000e-07 V_hig
+ 5.792000000e-07 V_hig
+ 5.792010000e-07 V_hig
+ 5.793000000e-07 V_hig
+ 5.793010000e-07 V_hig
+ 5.794000000e-07 V_hig
+ 5.794010000e-07 V_hig
+ 5.795000000e-07 V_hig
+ 5.795010000e-07 V_hig
+ 5.796000000e-07 V_hig
+ 5.796010000e-07 V_hig
+ 5.797000000e-07 V_hig
+ 5.797010000e-07 V_hig
+ 5.798000000e-07 V_hig
+ 5.798010000e-07 V_hig
+ 5.799000000e-07 V_hig
+ 5.799010000e-07 V_low
+ 5.800000000e-07 V_low
+ 5.800010000e-07 V_low
+ 5.801000000e-07 V_low
+ 5.801010000e-07 V_low
+ 5.802000000e-07 V_low
+ 5.802010000e-07 V_low
+ 5.803000000e-07 V_low
+ 5.803010000e-07 V_low
+ 5.804000000e-07 V_low
+ 5.804010000e-07 V_low
+ 5.805000000e-07 V_low
+ 5.805010000e-07 V_low
+ 5.806000000e-07 V_low
+ 5.806010000e-07 V_low
+ 5.807000000e-07 V_low
+ 5.807010000e-07 V_low
+ 5.808000000e-07 V_low
+ 5.808010000e-07 V_low
+ 5.809000000e-07 V_low
+ 5.809010000e-07 V_low
+ 5.810000000e-07 V_low
+ 5.810010000e-07 V_low
+ 5.811000000e-07 V_low
+ 5.811010000e-07 V_low
+ 5.812000000e-07 V_low
+ 5.812010000e-07 V_low
+ 5.813000000e-07 V_low
+ 5.813010000e-07 V_low
+ 5.814000000e-07 V_low
+ 5.814010000e-07 V_low
+ 5.815000000e-07 V_low
+ 5.815010000e-07 V_low
+ 5.816000000e-07 V_low
+ 5.816010000e-07 V_low
+ 5.817000000e-07 V_low
+ 5.817010000e-07 V_low
+ 5.818000000e-07 V_low
+ 5.818010000e-07 V_low
+ 5.819000000e-07 V_low
+ 5.819010000e-07 V_low
+ 5.820000000e-07 V_low
+ 5.820010000e-07 V_low
+ 5.821000000e-07 V_low
+ 5.821010000e-07 V_low
+ 5.822000000e-07 V_low
+ 5.822010000e-07 V_low
+ 5.823000000e-07 V_low
+ 5.823010000e-07 V_low
+ 5.824000000e-07 V_low
+ 5.824010000e-07 V_low
+ 5.825000000e-07 V_low
+ 5.825010000e-07 V_low
+ 5.826000000e-07 V_low
+ 5.826010000e-07 V_low
+ 5.827000000e-07 V_low
+ 5.827010000e-07 V_low
+ 5.828000000e-07 V_low
+ 5.828010000e-07 V_low
+ 5.829000000e-07 V_low
+ 5.829010000e-07 V_low
+ 5.830000000e-07 V_low
+ 5.830010000e-07 V_low
+ 5.831000000e-07 V_low
+ 5.831010000e-07 V_low
+ 5.832000000e-07 V_low
+ 5.832010000e-07 V_low
+ 5.833000000e-07 V_low
+ 5.833010000e-07 V_low
+ 5.834000000e-07 V_low
+ 5.834010000e-07 V_low
+ 5.835000000e-07 V_low
+ 5.835010000e-07 V_low
+ 5.836000000e-07 V_low
+ 5.836010000e-07 V_low
+ 5.837000000e-07 V_low
+ 5.837010000e-07 V_low
+ 5.838000000e-07 V_low
+ 5.838010000e-07 V_low
+ 5.839000000e-07 V_low
+ 5.839010000e-07 V_hig
+ 5.840000000e-07 V_hig
+ 5.840010000e-07 V_hig
+ 5.841000000e-07 V_hig
+ 5.841010000e-07 V_hig
+ 5.842000000e-07 V_hig
+ 5.842010000e-07 V_hig
+ 5.843000000e-07 V_hig
+ 5.843010000e-07 V_hig
+ 5.844000000e-07 V_hig
+ 5.844010000e-07 V_hig
+ 5.845000000e-07 V_hig
+ 5.845010000e-07 V_hig
+ 5.846000000e-07 V_hig
+ 5.846010000e-07 V_hig
+ 5.847000000e-07 V_hig
+ 5.847010000e-07 V_hig
+ 5.848000000e-07 V_hig
+ 5.848010000e-07 V_hig
+ 5.849000000e-07 V_hig
+ 5.849010000e-07 V_low
+ 5.850000000e-07 V_low
+ 5.850010000e-07 V_low
+ 5.851000000e-07 V_low
+ 5.851010000e-07 V_low
+ 5.852000000e-07 V_low
+ 5.852010000e-07 V_low
+ 5.853000000e-07 V_low
+ 5.853010000e-07 V_low
+ 5.854000000e-07 V_low
+ 5.854010000e-07 V_low
+ 5.855000000e-07 V_low
+ 5.855010000e-07 V_low
+ 5.856000000e-07 V_low
+ 5.856010000e-07 V_low
+ 5.857000000e-07 V_low
+ 5.857010000e-07 V_low
+ 5.858000000e-07 V_low
+ 5.858010000e-07 V_low
+ 5.859000000e-07 V_low
+ 5.859010000e-07 V_hig
+ 5.860000000e-07 V_hig
+ 5.860010000e-07 V_hig
+ 5.861000000e-07 V_hig
+ 5.861010000e-07 V_hig
+ 5.862000000e-07 V_hig
+ 5.862010000e-07 V_hig
+ 5.863000000e-07 V_hig
+ 5.863010000e-07 V_hig
+ 5.864000000e-07 V_hig
+ 5.864010000e-07 V_hig
+ 5.865000000e-07 V_hig
+ 5.865010000e-07 V_hig
+ 5.866000000e-07 V_hig
+ 5.866010000e-07 V_hig
+ 5.867000000e-07 V_hig
+ 5.867010000e-07 V_hig
+ 5.868000000e-07 V_hig
+ 5.868010000e-07 V_hig
+ 5.869000000e-07 V_hig
+ 5.869010000e-07 V_hig
+ 5.870000000e-07 V_hig
+ 5.870010000e-07 V_hig
+ 5.871000000e-07 V_hig
+ 5.871010000e-07 V_hig
+ 5.872000000e-07 V_hig
+ 5.872010000e-07 V_hig
+ 5.873000000e-07 V_hig
+ 5.873010000e-07 V_hig
+ 5.874000000e-07 V_hig
+ 5.874010000e-07 V_hig
+ 5.875000000e-07 V_hig
+ 5.875010000e-07 V_hig
+ 5.876000000e-07 V_hig
+ 5.876010000e-07 V_hig
+ 5.877000000e-07 V_hig
+ 5.877010000e-07 V_hig
+ 5.878000000e-07 V_hig
+ 5.878010000e-07 V_hig
+ 5.879000000e-07 V_hig
+ 5.879010000e-07 V_hig
+ 5.880000000e-07 V_hig
+ 5.880010000e-07 V_hig
+ 5.881000000e-07 V_hig
+ 5.881010000e-07 V_hig
+ 5.882000000e-07 V_hig
+ 5.882010000e-07 V_hig
+ 5.883000000e-07 V_hig
+ 5.883010000e-07 V_hig
+ 5.884000000e-07 V_hig
+ 5.884010000e-07 V_hig
+ 5.885000000e-07 V_hig
+ 5.885010000e-07 V_hig
+ 5.886000000e-07 V_hig
+ 5.886010000e-07 V_hig
+ 5.887000000e-07 V_hig
+ 5.887010000e-07 V_hig
+ 5.888000000e-07 V_hig
+ 5.888010000e-07 V_hig
+ 5.889000000e-07 V_hig
+ 5.889010000e-07 V_low
+ 5.890000000e-07 V_low
+ 5.890010000e-07 V_low
+ 5.891000000e-07 V_low
+ 5.891010000e-07 V_low
+ 5.892000000e-07 V_low
+ 5.892010000e-07 V_low
+ 5.893000000e-07 V_low
+ 5.893010000e-07 V_low
+ 5.894000000e-07 V_low
+ 5.894010000e-07 V_low
+ 5.895000000e-07 V_low
+ 5.895010000e-07 V_low
+ 5.896000000e-07 V_low
+ 5.896010000e-07 V_low
+ 5.897000000e-07 V_low
+ 5.897010000e-07 V_low
+ 5.898000000e-07 V_low
+ 5.898010000e-07 V_low
+ 5.899000000e-07 V_low
+ 5.899010000e-07 V_hig
+ 5.900000000e-07 V_hig
+ 5.900010000e-07 V_hig
+ 5.901000000e-07 V_hig
+ 5.901010000e-07 V_hig
+ 5.902000000e-07 V_hig
+ 5.902010000e-07 V_hig
+ 5.903000000e-07 V_hig
+ 5.903010000e-07 V_hig
+ 5.904000000e-07 V_hig
+ 5.904010000e-07 V_hig
+ 5.905000000e-07 V_hig
+ 5.905010000e-07 V_hig
+ 5.906000000e-07 V_hig
+ 5.906010000e-07 V_hig
+ 5.907000000e-07 V_hig
+ 5.907010000e-07 V_hig
+ 5.908000000e-07 V_hig
+ 5.908010000e-07 V_hig
+ 5.909000000e-07 V_hig
+ 5.909010000e-07 V_low
+ 5.910000000e-07 V_low
+ 5.910010000e-07 V_low
+ 5.911000000e-07 V_low
+ 5.911010000e-07 V_low
+ 5.912000000e-07 V_low
+ 5.912010000e-07 V_low
+ 5.913000000e-07 V_low
+ 5.913010000e-07 V_low
+ 5.914000000e-07 V_low
+ 5.914010000e-07 V_low
+ 5.915000000e-07 V_low
+ 5.915010000e-07 V_low
+ 5.916000000e-07 V_low
+ 5.916010000e-07 V_low
+ 5.917000000e-07 V_low
+ 5.917010000e-07 V_low
+ 5.918000000e-07 V_low
+ 5.918010000e-07 V_low
+ 5.919000000e-07 V_low
+ 5.919010000e-07 V_hig
+ 5.920000000e-07 V_hig
+ 5.920010000e-07 V_hig
+ 5.921000000e-07 V_hig
+ 5.921010000e-07 V_hig
+ 5.922000000e-07 V_hig
+ 5.922010000e-07 V_hig
+ 5.923000000e-07 V_hig
+ 5.923010000e-07 V_hig
+ 5.924000000e-07 V_hig
+ 5.924010000e-07 V_hig
+ 5.925000000e-07 V_hig
+ 5.925010000e-07 V_hig
+ 5.926000000e-07 V_hig
+ 5.926010000e-07 V_hig
+ 5.927000000e-07 V_hig
+ 5.927010000e-07 V_hig
+ 5.928000000e-07 V_hig
+ 5.928010000e-07 V_hig
+ 5.929000000e-07 V_hig
+ 5.929010000e-07 V_hig
+ 5.930000000e-07 V_hig
+ 5.930010000e-07 V_hig
+ 5.931000000e-07 V_hig
+ 5.931010000e-07 V_hig
+ 5.932000000e-07 V_hig
+ 5.932010000e-07 V_hig
+ 5.933000000e-07 V_hig
+ 5.933010000e-07 V_hig
+ 5.934000000e-07 V_hig
+ 5.934010000e-07 V_hig
+ 5.935000000e-07 V_hig
+ 5.935010000e-07 V_hig
+ 5.936000000e-07 V_hig
+ 5.936010000e-07 V_hig
+ 5.937000000e-07 V_hig
+ 5.937010000e-07 V_hig
+ 5.938000000e-07 V_hig
+ 5.938010000e-07 V_hig
+ 5.939000000e-07 V_hig
+ 5.939010000e-07 V_hig
+ 5.940000000e-07 V_hig
+ 5.940010000e-07 V_hig
+ 5.941000000e-07 V_hig
+ 5.941010000e-07 V_hig
+ 5.942000000e-07 V_hig
+ 5.942010000e-07 V_hig
+ 5.943000000e-07 V_hig
+ 5.943010000e-07 V_hig
+ 5.944000000e-07 V_hig
+ 5.944010000e-07 V_hig
+ 5.945000000e-07 V_hig
+ 5.945010000e-07 V_hig
+ 5.946000000e-07 V_hig
+ 5.946010000e-07 V_hig
+ 5.947000000e-07 V_hig
+ 5.947010000e-07 V_hig
+ 5.948000000e-07 V_hig
+ 5.948010000e-07 V_hig
+ 5.949000000e-07 V_hig
+ 5.949010000e-07 V_hig
+ 5.950000000e-07 V_hig
+ 5.950010000e-07 V_hig
+ 5.951000000e-07 V_hig
+ 5.951010000e-07 V_hig
+ 5.952000000e-07 V_hig
+ 5.952010000e-07 V_hig
+ 5.953000000e-07 V_hig
+ 5.953010000e-07 V_hig
+ 5.954000000e-07 V_hig
+ 5.954010000e-07 V_hig
+ 5.955000000e-07 V_hig
+ 5.955010000e-07 V_hig
+ 5.956000000e-07 V_hig
+ 5.956010000e-07 V_hig
+ 5.957000000e-07 V_hig
+ 5.957010000e-07 V_hig
+ 5.958000000e-07 V_hig
+ 5.958010000e-07 V_hig
+ 5.959000000e-07 V_hig
+ 5.959010000e-07 V_hig
+ 5.960000000e-07 V_hig
+ 5.960010000e-07 V_hig
+ 5.961000000e-07 V_hig
+ 5.961010000e-07 V_hig
+ 5.962000000e-07 V_hig
+ 5.962010000e-07 V_hig
+ 5.963000000e-07 V_hig
+ 5.963010000e-07 V_hig
+ 5.964000000e-07 V_hig
+ 5.964010000e-07 V_hig
+ 5.965000000e-07 V_hig
+ 5.965010000e-07 V_hig
+ 5.966000000e-07 V_hig
+ 5.966010000e-07 V_hig
+ 5.967000000e-07 V_hig
+ 5.967010000e-07 V_hig
+ 5.968000000e-07 V_hig
+ 5.968010000e-07 V_hig
+ 5.969000000e-07 V_hig
+ 5.969010000e-07 V_low
+ 5.970000000e-07 V_low
+ 5.970010000e-07 V_low
+ 5.971000000e-07 V_low
+ 5.971010000e-07 V_low
+ 5.972000000e-07 V_low
+ 5.972010000e-07 V_low
+ 5.973000000e-07 V_low
+ 5.973010000e-07 V_low
+ 5.974000000e-07 V_low
+ 5.974010000e-07 V_low
+ 5.975000000e-07 V_low
+ 5.975010000e-07 V_low
+ 5.976000000e-07 V_low
+ 5.976010000e-07 V_low
+ 5.977000000e-07 V_low
+ 5.977010000e-07 V_low
+ 5.978000000e-07 V_low
+ 5.978010000e-07 V_low
+ 5.979000000e-07 V_low
+ 5.979010000e-07 V_hig
+ 5.980000000e-07 V_hig
+ 5.980010000e-07 V_hig
+ 5.981000000e-07 V_hig
+ 5.981010000e-07 V_hig
+ 5.982000000e-07 V_hig
+ 5.982010000e-07 V_hig
+ 5.983000000e-07 V_hig
+ 5.983010000e-07 V_hig
+ 5.984000000e-07 V_hig
+ 5.984010000e-07 V_hig
+ 5.985000000e-07 V_hig
+ 5.985010000e-07 V_hig
+ 5.986000000e-07 V_hig
+ 5.986010000e-07 V_hig
+ 5.987000000e-07 V_hig
+ 5.987010000e-07 V_hig
+ 5.988000000e-07 V_hig
+ 5.988010000e-07 V_hig
+ 5.989000000e-07 V_hig
+ 5.989010000e-07 V_hig
+ 5.990000000e-07 V_hig
+ 5.990010000e-07 V_hig
+ 5.991000000e-07 V_hig
+ 5.991010000e-07 V_hig
+ 5.992000000e-07 V_hig
+ 5.992010000e-07 V_hig
+ 5.993000000e-07 V_hig
+ 5.993010000e-07 V_hig
+ 5.994000000e-07 V_hig
+ 5.994010000e-07 V_hig
+ 5.995000000e-07 V_hig
+ 5.995010000e-07 V_hig
+ 5.996000000e-07 V_hig
+ 5.996010000e-07 V_hig
+ 5.997000000e-07 V_hig
+ 5.997010000e-07 V_hig
+ 5.998000000e-07 V_hig
+ 5.998010000e-07 V_hig
+ 5.999000000e-07 V_hig
+ 5.999010000e-07 V_hig
+ 6.000000000e-07 V_hig
+ 6.000010000e-07 V_hig
+ 6.001000000e-07 V_hig
+ 6.001010000e-07 V_hig
+ 6.002000000e-07 V_hig
+ 6.002010000e-07 V_hig
+ 6.003000000e-07 V_hig
+ 6.003010000e-07 V_hig
+ 6.004000000e-07 V_hig
+ 6.004010000e-07 V_hig
+ 6.005000000e-07 V_hig
+ 6.005010000e-07 V_hig
+ 6.006000000e-07 V_hig
+ 6.006010000e-07 V_hig
+ 6.007000000e-07 V_hig
+ 6.007010000e-07 V_hig
+ 6.008000000e-07 V_hig
+ 6.008010000e-07 V_hig
+ 6.009000000e-07 V_hig
+ 6.009010000e-07 V_low
+ 6.010000000e-07 V_low
+ 6.010010000e-07 V_low
+ 6.011000000e-07 V_low
+ 6.011010000e-07 V_low
+ 6.012000000e-07 V_low
+ 6.012010000e-07 V_low
+ 6.013000000e-07 V_low
+ 6.013010000e-07 V_low
+ 6.014000000e-07 V_low
+ 6.014010000e-07 V_low
+ 6.015000000e-07 V_low
+ 6.015010000e-07 V_low
+ 6.016000000e-07 V_low
+ 6.016010000e-07 V_low
+ 6.017000000e-07 V_low
+ 6.017010000e-07 V_low
+ 6.018000000e-07 V_low
+ 6.018010000e-07 V_low
+ 6.019000000e-07 V_low
+ 6.019010000e-07 V_low
+ 6.020000000e-07 V_low
+ 6.020010000e-07 V_low
+ 6.021000000e-07 V_low
+ 6.021010000e-07 V_low
+ 6.022000000e-07 V_low
+ 6.022010000e-07 V_low
+ 6.023000000e-07 V_low
+ 6.023010000e-07 V_low
+ 6.024000000e-07 V_low
+ 6.024010000e-07 V_low
+ 6.025000000e-07 V_low
+ 6.025010000e-07 V_low
+ 6.026000000e-07 V_low
+ 6.026010000e-07 V_low
+ 6.027000000e-07 V_low
+ 6.027010000e-07 V_low
+ 6.028000000e-07 V_low
+ 6.028010000e-07 V_low
+ 6.029000000e-07 V_low
+ 6.029010000e-07 V_low
+ 6.030000000e-07 V_low
+ 6.030010000e-07 V_low
+ 6.031000000e-07 V_low
+ 6.031010000e-07 V_low
+ 6.032000000e-07 V_low
+ 6.032010000e-07 V_low
+ 6.033000000e-07 V_low
+ 6.033010000e-07 V_low
+ 6.034000000e-07 V_low
+ 6.034010000e-07 V_low
+ 6.035000000e-07 V_low
+ 6.035010000e-07 V_low
+ 6.036000000e-07 V_low
+ 6.036010000e-07 V_low
+ 6.037000000e-07 V_low
+ 6.037010000e-07 V_low
+ 6.038000000e-07 V_low
+ 6.038010000e-07 V_low
+ 6.039000000e-07 V_low
+ 6.039010000e-07 V_hig
+ 6.040000000e-07 V_hig
+ 6.040010000e-07 V_hig
+ 6.041000000e-07 V_hig
+ 6.041010000e-07 V_hig
+ 6.042000000e-07 V_hig
+ 6.042010000e-07 V_hig
+ 6.043000000e-07 V_hig
+ 6.043010000e-07 V_hig
+ 6.044000000e-07 V_hig
+ 6.044010000e-07 V_hig
+ 6.045000000e-07 V_hig
+ 6.045010000e-07 V_hig
+ 6.046000000e-07 V_hig
+ 6.046010000e-07 V_hig
+ 6.047000000e-07 V_hig
+ 6.047010000e-07 V_hig
+ 6.048000000e-07 V_hig
+ 6.048010000e-07 V_hig
+ 6.049000000e-07 V_hig
+ 6.049010000e-07 V_hig
+ 6.050000000e-07 V_hig
+ 6.050010000e-07 V_hig
+ 6.051000000e-07 V_hig
+ 6.051010000e-07 V_hig
+ 6.052000000e-07 V_hig
+ 6.052010000e-07 V_hig
+ 6.053000000e-07 V_hig
+ 6.053010000e-07 V_hig
+ 6.054000000e-07 V_hig
+ 6.054010000e-07 V_hig
+ 6.055000000e-07 V_hig
+ 6.055010000e-07 V_hig
+ 6.056000000e-07 V_hig
+ 6.056010000e-07 V_hig
+ 6.057000000e-07 V_hig
+ 6.057010000e-07 V_hig
+ 6.058000000e-07 V_hig
+ 6.058010000e-07 V_hig
+ 6.059000000e-07 V_hig
+ 6.059010000e-07 V_hig
+ 6.060000000e-07 V_hig
+ 6.060010000e-07 V_hig
+ 6.061000000e-07 V_hig
+ 6.061010000e-07 V_hig
+ 6.062000000e-07 V_hig
+ 6.062010000e-07 V_hig
+ 6.063000000e-07 V_hig
+ 6.063010000e-07 V_hig
+ 6.064000000e-07 V_hig
+ 6.064010000e-07 V_hig
+ 6.065000000e-07 V_hig
+ 6.065010000e-07 V_hig
+ 6.066000000e-07 V_hig
+ 6.066010000e-07 V_hig
+ 6.067000000e-07 V_hig
+ 6.067010000e-07 V_hig
+ 6.068000000e-07 V_hig
+ 6.068010000e-07 V_hig
+ 6.069000000e-07 V_hig
+ 6.069010000e-07 V_hig
+ 6.070000000e-07 V_hig
+ 6.070010000e-07 V_hig
+ 6.071000000e-07 V_hig
+ 6.071010000e-07 V_hig
+ 6.072000000e-07 V_hig
+ 6.072010000e-07 V_hig
+ 6.073000000e-07 V_hig
+ 6.073010000e-07 V_hig
+ 6.074000000e-07 V_hig
+ 6.074010000e-07 V_hig
+ 6.075000000e-07 V_hig
+ 6.075010000e-07 V_hig
+ 6.076000000e-07 V_hig
+ 6.076010000e-07 V_hig
+ 6.077000000e-07 V_hig
+ 6.077010000e-07 V_hig
+ 6.078000000e-07 V_hig
+ 6.078010000e-07 V_hig
+ 6.079000000e-07 V_hig
+ 6.079010000e-07 V_hig
+ 6.080000000e-07 V_hig
+ 6.080010000e-07 V_hig
+ 6.081000000e-07 V_hig
+ 6.081010000e-07 V_hig
+ 6.082000000e-07 V_hig
+ 6.082010000e-07 V_hig
+ 6.083000000e-07 V_hig
+ 6.083010000e-07 V_hig
+ 6.084000000e-07 V_hig
+ 6.084010000e-07 V_hig
+ 6.085000000e-07 V_hig
+ 6.085010000e-07 V_hig
+ 6.086000000e-07 V_hig
+ 6.086010000e-07 V_hig
+ 6.087000000e-07 V_hig
+ 6.087010000e-07 V_hig
+ 6.088000000e-07 V_hig
+ 6.088010000e-07 V_hig
+ 6.089000000e-07 V_hig
+ 6.089010000e-07 V_low
+ 6.090000000e-07 V_low
+ 6.090010000e-07 V_low
+ 6.091000000e-07 V_low
+ 6.091010000e-07 V_low
+ 6.092000000e-07 V_low
+ 6.092010000e-07 V_low
+ 6.093000000e-07 V_low
+ 6.093010000e-07 V_low
+ 6.094000000e-07 V_low
+ 6.094010000e-07 V_low
+ 6.095000000e-07 V_low
+ 6.095010000e-07 V_low
+ 6.096000000e-07 V_low
+ 6.096010000e-07 V_low
+ 6.097000000e-07 V_low
+ 6.097010000e-07 V_low
+ 6.098000000e-07 V_low
+ 6.098010000e-07 V_low
+ 6.099000000e-07 V_low
+ 6.099010000e-07 V_low
+ 6.100000000e-07 V_low
+ 6.100010000e-07 V_low
+ 6.101000000e-07 V_low
+ 6.101010000e-07 V_low
+ 6.102000000e-07 V_low
+ 6.102010000e-07 V_low
+ 6.103000000e-07 V_low
+ 6.103010000e-07 V_low
+ 6.104000000e-07 V_low
+ 6.104010000e-07 V_low
+ 6.105000000e-07 V_low
+ 6.105010000e-07 V_low
+ 6.106000000e-07 V_low
+ 6.106010000e-07 V_low
+ 6.107000000e-07 V_low
+ 6.107010000e-07 V_low
+ 6.108000000e-07 V_low
+ 6.108010000e-07 V_low
+ 6.109000000e-07 V_low
+ 6.109010000e-07 V_hig
+ 6.110000000e-07 V_hig
+ 6.110010000e-07 V_hig
+ 6.111000000e-07 V_hig
+ 6.111010000e-07 V_hig
+ 6.112000000e-07 V_hig
+ 6.112010000e-07 V_hig
+ 6.113000000e-07 V_hig
+ 6.113010000e-07 V_hig
+ 6.114000000e-07 V_hig
+ 6.114010000e-07 V_hig
+ 6.115000000e-07 V_hig
+ 6.115010000e-07 V_hig
+ 6.116000000e-07 V_hig
+ 6.116010000e-07 V_hig
+ 6.117000000e-07 V_hig
+ 6.117010000e-07 V_hig
+ 6.118000000e-07 V_hig
+ 6.118010000e-07 V_hig
+ 6.119000000e-07 V_hig
+ 6.119010000e-07 V_low
+ 6.120000000e-07 V_low
+ 6.120010000e-07 V_low
+ 6.121000000e-07 V_low
+ 6.121010000e-07 V_low
+ 6.122000000e-07 V_low
+ 6.122010000e-07 V_low
+ 6.123000000e-07 V_low
+ 6.123010000e-07 V_low
+ 6.124000000e-07 V_low
+ 6.124010000e-07 V_low
+ 6.125000000e-07 V_low
+ 6.125010000e-07 V_low
+ 6.126000000e-07 V_low
+ 6.126010000e-07 V_low
+ 6.127000000e-07 V_low
+ 6.127010000e-07 V_low
+ 6.128000000e-07 V_low
+ 6.128010000e-07 V_low
+ 6.129000000e-07 V_low
+ 6.129010000e-07 V_hig
+ 6.130000000e-07 V_hig
+ 6.130010000e-07 V_hig
+ 6.131000000e-07 V_hig
+ 6.131010000e-07 V_hig
+ 6.132000000e-07 V_hig
+ 6.132010000e-07 V_hig
+ 6.133000000e-07 V_hig
+ 6.133010000e-07 V_hig
+ 6.134000000e-07 V_hig
+ 6.134010000e-07 V_hig
+ 6.135000000e-07 V_hig
+ 6.135010000e-07 V_hig
+ 6.136000000e-07 V_hig
+ 6.136010000e-07 V_hig
+ 6.137000000e-07 V_hig
+ 6.137010000e-07 V_hig
+ 6.138000000e-07 V_hig
+ 6.138010000e-07 V_hig
+ 6.139000000e-07 V_hig
+ 6.139010000e-07 V_hig
+ 6.140000000e-07 V_hig
+ 6.140010000e-07 V_hig
+ 6.141000000e-07 V_hig
+ 6.141010000e-07 V_hig
+ 6.142000000e-07 V_hig
+ 6.142010000e-07 V_hig
+ 6.143000000e-07 V_hig
+ 6.143010000e-07 V_hig
+ 6.144000000e-07 V_hig
+ 6.144010000e-07 V_hig
+ 6.145000000e-07 V_hig
+ 6.145010000e-07 V_hig
+ 6.146000000e-07 V_hig
+ 6.146010000e-07 V_hig
+ 6.147000000e-07 V_hig
+ 6.147010000e-07 V_hig
+ 6.148000000e-07 V_hig
+ 6.148010000e-07 V_hig
+ 6.149000000e-07 V_hig
+ 6.149010000e-07 V_hig
+ 6.150000000e-07 V_hig
+ 6.150010000e-07 V_hig
+ 6.151000000e-07 V_hig
+ 6.151010000e-07 V_hig
+ 6.152000000e-07 V_hig
+ 6.152010000e-07 V_hig
+ 6.153000000e-07 V_hig
+ 6.153010000e-07 V_hig
+ 6.154000000e-07 V_hig
+ 6.154010000e-07 V_hig
+ 6.155000000e-07 V_hig
+ 6.155010000e-07 V_hig
+ 6.156000000e-07 V_hig
+ 6.156010000e-07 V_hig
+ 6.157000000e-07 V_hig
+ 6.157010000e-07 V_hig
+ 6.158000000e-07 V_hig
+ 6.158010000e-07 V_hig
+ 6.159000000e-07 V_hig
+ 6.159010000e-07 V_hig
+ 6.160000000e-07 V_hig
+ 6.160010000e-07 V_hig
+ 6.161000000e-07 V_hig
+ 6.161010000e-07 V_hig
+ 6.162000000e-07 V_hig
+ 6.162010000e-07 V_hig
+ 6.163000000e-07 V_hig
+ 6.163010000e-07 V_hig
+ 6.164000000e-07 V_hig
+ 6.164010000e-07 V_hig
+ 6.165000000e-07 V_hig
+ 6.165010000e-07 V_hig
+ 6.166000000e-07 V_hig
+ 6.166010000e-07 V_hig
+ 6.167000000e-07 V_hig
+ 6.167010000e-07 V_hig
+ 6.168000000e-07 V_hig
+ 6.168010000e-07 V_hig
+ 6.169000000e-07 V_hig
+ 6.169010000e-07 V_hig
+ 6.170000000e-07 V_hig
+ 6.170010000e-07 V_hig
+ 6.171000000e-07 V_hig
+ 6.171010000e-07 V_hig
+ 6.172000000e-07 V_hig
+ 6.172010000e-07 V_hig
+ 6.173000000e-07 V_hig
+ 6.173010000e-07 V_hig
+ 6.174000000e-07 V_hig
+ 6.174010000e-07 V_hig
+ 6.175000000e-07 V_hig
+ 6.175010000e-07 V_hig
+ 6.176000000e-07 V_hig
+ 6.176010000e-07 V_hig
+ 6.177000000e-07 V_hig
+ 6.177010000e-07 V_hig
+ 6.178000000e-07 V_hig
+ 6.178010000e-07 V_hig
+ 6.179000000e-07 V_hig
+ 6.179010000e-07 V_hig
+ 6.180000000e-07 V_hig
+ 6.180010000e-07 V_hig
+ 6.181000000e-07 V_hig
+ 6.181010000e-07 V_hig
+ 6.182000000e-07 V_hig
+ 6.182010000e-07 V_hig
+ 6.183000000e-07 V_hig
+ 6.183010000e-07 V_hig
+ 6.184000000e-07 V_hig
+ 6.184010000e-07 V_hig
+ 6.185000000e-07 V_hig
+ 6.185010000e-07 V_hig
+ 6.186000000e-07 V_hig
+ 6.186010000e-07 V_hig
+ 6.187000000e-07 V_hig
+ 6.187010000e-07 V_hig
+ 6.188000000e-07 V_hig
+ 6.188010000e-07 V_hig
+ 6.189000000e-07 V_hig
+ 6.189010000e-07 V_hig
+ 6.190000000e-07 V_hig
+ 6.190010000e-07 V_hig
+ 6.191000000e-07 V_hig
+ 6.191010000e-07 V_hig
+ 6.192000000e-07 V_hig
+ 6.192010000e-07 V_hig
+ 6.193000000e-07 V_hig
+ 6.193010000e-07 V_hig
+ 6.194000000e-07 V_hig
+ 6.194010000e-07 V_hig
+ 6.195000000e-07 V_hig
+ 6.195010000e-07 V_hig
+ 6.196000000e-07 V_hig
+ 6.196010000e-07 V_hig
+ 6.197000000e-07 V_hig
+ 6.197010000e-07 V_hig
+ 6.198000000e-07 V_hig
+ 6.198010000e-07 V_hig
+ 6.199000000e-07 V_hig
+ 6.199010000e-07 V_hig
+ 6.200000000e-07 V_hig
+ 6.200010000e-07 V_hig
+ 6.201000000e-07 V_hig
+ 6.201010000e-07 V_hig
+ 6.202000000e-07 V_hig
+ 6.202010000e-07 V_hig
+ 6.203000000e-07 V_hig
+ 6.203010000e-07 V_hig
+ 6.204000000e-07 V_hig
+ 6.204010000e-07 V_hig
+ 6.205000000e-07 V_hig
+ 6.205010000e-07 V_hig
+ 6.206000000e-07 V_hig
+ 6.206010000e-07 V_hig
+ 6.207000000e-07 V_hig
+ 6.207010000e-07 V_hig
+ 6.208000000e-07 V_hig
+ 6.208010000e-07 V_hig
+ 6.209000000e-07 V_hig
+ 6.209010000e-07 V_hig
+ 6.210000000e-07 V_hig
+ 6.210010000e-07 V_hig
+ 6.211000000e-07 V_hig
+ 6.211010000e-07 V_hig
+ 6.212000000e-07 V_hig
+ 6.212010000e-07 V_hig
+ 6.213000000e-07 V_hig
+ 6.213010000e-07 V_hig
+ 6.214000000e-07 V_hig
+ 6.214010000e-07 V_hig
+ 6.215000000e-07 V_hig
+ 6.215010000e-07 V_hig
+ 6.216000000e-07 V_hig
+ 6.216010000e-07 V_hig
+ 6.217000000e-07 V_hig
+ 6.217010000e-07 V_hig
+ 6.218000000e-07 V_hig
+ 6.218010000e-07 V_hig
+ 6.219000000e-07 V_hig
+ 6.219010000e-07 V_low
+ 6.220000000e-07 V_low
+ 6.220010000e-07 V_low
+ 6.221000000e-07 V_low
+ 6.221010000e-07 V_low
+ 6.222000000e-07 V_low
+ 6.222010000e-07 V_low
+ 6.223000000e-07 V_low
+ 6.223010000e-07 V_low
+ 6.224000000e-07 V_low
+ 6.224010000e-07 V_low
+ 6.225000000e-07 V_low
+ 6.225010000e-07 V_low
+ 6.226000000e-07 V_low
+ 6.226010000e-07 V_low
+ 6.227000000e-07 V_low
+ 6.227010000e-07 V_low
+ 6.228000000e-07 V_low
+ 6.228010000e-07 V_low
+ 6.229000000e-07 V_low
+ 6.229010000e-07 V_hig
+ 6.230000000e-07 V_hig
+ 6.230010000e-07 V_hig
+ 6.231000000e-07 V_hig
+ 6.231010000e-07 V_hig
+ 6.232000000e-07 V_hig
+ 6.232010000e-07 V_hig
+ 6.233000000e-07 V_hig
+ 6.233010000e-07 V_hig
+ 6.234000000e-07 V_hig
+ 6.234010000e-07 V_hig
+ 6.235000000e-07 V_hig
+ 6.235010000e-07 V_hig
+ 6.236000000e-07 V_hig
+ 6.236010000e-07 V_hig
+ 6.237000000e-07 V_hig
+ 6.237010000e-07 V_hig
+ 6.238000000e-07 V_hig
+ 6.238010000e-07 V_hig
+ 6.239000000e-07 V_hig
+ 6.239010000e-07 V_low
+ 6.240000000e-07 V_low
+ 6.240010000e-07 V_low
+ 6.241000000e-07 V_low
+ 6.241010000e-07 V_low
+ 6.242000000e-07 V_low
+ 6.242010000e-07 V_low
+ 6.243000000e-07 V_low
+ 6.243010000e-07 V_low
+ 6.244000000e-07 V_low
+ 6.244010000e-07 V_low
+ 6.245000000e-07 V_low
+ 6.245010000e-07 V_low
+ 6.246000000e-07 V_low
+ 6.246010000e-07 V_low
+ 6.247000000e-07 V_low
+ 6.247010000e-07 V_low
+ 6.248000000e-07 V_low
+ 6.248010000e-07 V_low
+ 6.249000000e-07 V_low
+ 6.249010000e-07 V_hig
+ 6.250000000e-07 V_hig
+ 6.250010000e-07 V_hig
+ 6.251000000e-07 V_hig
+ 6.251010000e-07 V_hig
+ 6.252000000e-07 V_hig
+ 6.252010000e-07 V_hig
+ 6.253000000e-07 V_hig
+ 6.253010000e-07 V_hig
+ 6.254000000e-07 V_hig
+ 6.254010000e-07 V_hig
+ 6.255000000e-07 V_hig
+ 6.255010000e-07 V_hig
+ 6.256000000e-07 V_hig
+ 6.256010000e-07 V_hig
+ 6.257000000e-07 V_hig
+ 6.257010000e-07 V_hig
+ 6.258000000e-07 V_hig
+ 6.258010000e-07 V_hig
+ 6.259000000e-07 V_hig
+ 6.259010000e-07 V_low
+ 6.260000000e-07 V_low
+ 6.260010000e-07 V_low
+ 6.261000000e-07 V_low
+ 6.261010000e-07 V_low
+ 6.262000000e-07 V_low
+ 6.262010000e-07 V_low
+ 6.263000000e-07 V_low
+ 6.263010000e-07 V_low
+ 6.264000000e-07 V_low
+ 6.264010000e-07 V_low
+ 6.265000000e-07 V_low
+ 6.265010000e-07 V_low
+ 6.266000000e-07 V_low
+ 6.266010000e-07 V_low
+ 6.267000000e-07 V_low
+ 6.267010000e-07 V_low
+ 6.268000000e-07 V_low
+ 6.268010000e-07 V_low
+ 6.269000000e-07 V_low
+ 6.269010000e-07 V_low
+ 6.270000000e-07 V_low
+ 6.270010000e-07 V_low
+ 6.271000000e-07 V_low
+ 6.271010000e-07 V_low
+ 6.272000000e-07 V_low
+ 6.272010000e-07 V_low
+ 6.273000000e-07 V_low
+ 6.273010000e-07 V_low
+ 6.274000000e-07 V_low
+ 6.274010000e-07 V_low
+ 6.275000000e-07 V_low
+ 6.275010000e-07 V_low
+ 6.276000000e-07 V_low
+ 6.276010000e-07 V_low
+ 6.277000000e-07 V_low
+ 6.277010000e-07 V_low
+ 6.278000000e-07 V_low
+ 6.278010000e-07 V_low
+ 6.279000000e-07 V_low
+ 6.279010000e-07 V_hig
+ 6.280000000e-07 V_hig
+ 6.280010000e-07 V_hig
+ 6.281000000e-07 V_hig
+ 6.281010000e-07 V_hig
+ 6.282000000e-07 V_hig
+ 6.282010000e-07 V_hig
+ 6.283000000e-07 V_hig
+ 6.283010000e-07 V_hig
+ 6.284000000e-07 V_hig
+ 6.284010000e-07 V_hig
+ 6.285000000e-07 V_hig
+ 6.285010000e-07 V_hig
+ 6.286000000e-07 V_hig
+ 6.286010000e-07 V_hig
+ 6.287000000e-07 V_hig
+ 6.287010000e-07 V_hig
+ 6.288000000e-07 V_hig
+ 6.288010000e-07 V_hig
+ 6.289000000e-07 V_hig
+ 6.289010000e-07 V_hig
+ 6.290000000e-07 V_hig
+ 6.290010000e-07 V_hig
+ 6.291000000e-07 V_hig
+ 6.291010000e-07 V_hig
+ 6.292000000e-07 V_hig
+ 6.292010000e-07 V_hig
+ 6.293000000e-07 V_hig
+ 6.293010000e-07 V_hig
+ 6.294000000e-07 V_hig
+ 6.294010000e-07 V_hig
+ 6.295000000e-07 V_hig
+ 6.295010000e-07 V_hig
+ 6.296000000e-07 V_hig
+ 6.296010000e-07 V_hig
+ 6.297000000e-07 V_hig
+ 6.297010000e-07 V_hig
+ 6.298000000e-07 V_hig
+ 6.298010000e-07 V_hig
+ 6.299000000e-07 V_hig
+ 6.299010000e-07 V_low
+ 6.300000000e-07 V_low
+ 6.300010000e-07 V_low
+ 6.301000000e-07 V_low
+ 6.301010000e-07 V_low
+ 6.302000000e-07 V_low
+ 6.302010000e-07 V_low
+ 6.303000000e-07 V_low
+ 6.303010000e-07 V_low
+ 6.304000000e-07 V_low
+ 6.304010000e-07 V_low
+ 6.305000000e-07 V_low
+ 6.305010000e-07 V_low
+ 6.306000000e-07 V_low
+ 6.306010000e-07 V_low
+ 6.307000000e-07 V_low
+ 6.307010000e-07 V_low
+ 6.308000000e-07 V_low
+ 6.308010000e-07 V_low
+ 6.309000000e-07 V_low
+ 6.309010000e-07 V_low
+ 6.310000000e-07 V_low
+ 6.310010000e-07 V_low
+ 6.311000000e-07 V_low
+ 6.311010000e-07 V_low
+ 6.312000000e-07 V_low
+ 6.312010000e-07 V_low
+ 6.313000000e-07 V_low
+ 6.313010000e-07 V_low
+ 6.314000000e-07 V_low
+ 6.314010000e-07 V_low
+ 6.315000000e-07 V_low
+ 6.315010000e-07 V_low
+ 6.316000000e-07 V_low
+ 6.316010000e-07 V_low
+ 6.317000000e-07 V_low
+ 6.317010000e-07 V_low
+ 6.318000000e-07 V_low
+ 6.318010000e-07 V_low
+ 6.319000000e-07 V_low
+ 6.319010000e-07 V_low
+ 6.320000000e-07 V_low
+ 6.320010000e-07 V_low
+ 6.321000000e-07 V_low
+ 6.321010000e-07 V_low
+ 6.322000000e-07 V_low
+ 6.322010000e-07 V_low
+ 6.323000000e-07 V_low
+ 6.323010000e-07 V_low
+ 6.324000000e-07 V_low
+ 6.324010000e-07 V_low
+ 6.325000000e-07 V_low
+ 6.325010000e-07 V_low
+ 6.326000000e-07 V_low
+ 6.326010000e-07 V_low
+ 6.327000000e-07 V_low
+ 6.327010000e-07 V_low
+ 6.328000000e-07 V_low
+ 6.328010000e-07 V_low
+ 6.329000000e-07 V_low
+ 6.329010000e-07 V_hig
+ 6.330000000e-07 V_hig
+ 6.330010000e-07 V_hig
+ 6.331000000e-07 V_hig
+ 6.331010000e-07 V_hig
+ 6.332000000e-07 V_hig
+ 6.332010000e-07 V_hig
+ 6.333000000e-07 V_hig
+ 6.333010000e-07 V_hig
+ 6.334000000e-07 V_hig
+ 6.334010000e-07 V_hig
+ 6.335000000e-07 V_hig
+ 6.335010000e-07 V_hig
+ 6.336000000e-07 V_hig
+ 6.336010000e-07 V_hig
+ 6.337000000e-07 V_hig
+ 6.337010000e-07 V_hig
+ 6.338000000e-07 V_hig
+ 6.338010000e-07 V_hig
+ 6.339000000e-07 V_hig
+ 6.339010000e-07 V_low
+ 6.340000000e-07 V_low
+ 6.340010000e-07 V_low
+ 6.341000000e-07 V_low
+ 6.341010000e-07 V_low
+ 6.342000000e-07 V_low
+ 6.342010000e-07 V_low
+ 6.343000000e-07 V_low
+ 6.343010000e-07 V_low
+ 6.344000000e-07 V_low
+ 6.344010000e-07 V_low
+ 6.345000000e-07 V_low
+ 6.345010000e-07 V_low
+ 6.346000000e-07 V_low
+ 6.346010000e-07 V_low
+ 6.347000000e-07 V_low
+ 6.347010000e-07 V_low
+ 6.348000000e-07 V_low
+ 6.348010000e-07 V_low
+ 6.349000000e-07 V_low
+ 6.349010000e-07 V_low
+ 6.350000000e-07 V_low
+ 6.350010000e-07 V_low
+ 6.351000000e-07 V_low
+ 6.351010000e-07 V_low
+ 6.352000000e-07 V_low
+ 6.352010000e-07 V_low
+ 6.353000000e-07 V_low
+ 6.353010000e-07 V_low
+ 6.354000000e-07 V_low
+ 6.354010000e-07 V_low
+ 6.355000000e-07 V_low
+ 6.355010000e-07 V_low
+ 6.356000000e-07 V_low
+ 6.356010000e-07 V_low
+ 6.357000000e-07 V_low
+ 6.357010000e-07 V_low
+ 6.358000000e-07 V_low
+ 6.358010000e-07 V_low
+ 6.359000000e-07 V_low
+ 6.359010000e-07 V_low
+ 6.360000000e-07 V_low
+ 6.360010000e-07 V_low
+ 6.361000000e-07 V_low
+ 6.361010000e-07 V_low
+ 6.362000000e-07 V_low
+ 6.362010000e-07 V_low
+ 6.363000000e-07 V_low
+ 6.363010000e-07 V_low
+ 6.364000000e-07 V_low
+ 6.364010000e-07 V_low
+ 6.365000000e-07 V_low
+ 6.365010000e-07 V_low
+ 6.366000000e-07 V_low
+ 6.366010000e-07 V_low
+ 6.367000000e-07 V_low
+ 6.367010000e-07 V_low
+ 6.368000000e-07 V_low
+ 6.368010000e-07 V_low
+ 6.369000000e-07 V_low
+ 6.369010000e-07 V_hig
+ 6.370000000e-07 V_hig
+ 6.370010000e-07 V_hig
+ 6.371000000e-07 V_hig
+ 6.371010000e-07 V_hig
+ 6.372000000e-07 V_hig
+ 6.372010000e-07 V_hig
+ 6.373000000e-07 V_hig
+ 6.373010000e-07 V_hig
+ 6.374000000e-07 V_hig
+ 6.374010000e-07 V_hig
+ 6.375000000e-07 V_hig
+ 6.375010000e-07 V_hig
+ 6.376000000e-07 V_hig
+ 6.376010000e-07 V_hig
+ 6.377000000e-07 V_hig
+ 6.377010000e-07 V_hig
+ 6.378000000e-07 V_hig
+ 6.378010000e-07 V_hig
+ 6.379000000e-07 V_hig
+ 6.379010000e-07 V_low
+ 6.380000000e-07 V_low
+ 6.380010000e-07 V_low
+ 6.381000000e-07 V_low
+ 6.381010000e-07 V_low
+ 6.382000000e-07 V_low
+ 6.382010000e-07 V_low
+ 6.383000000e-07 V_low
+ 6.383010000e-07 V_low
+ 6.384000000e-07 V_low
+ 6.384010000e-07 V_low
+ 6.385000000e-07 V_low
+ 6.385010000e-07 V_low
+ 6.386000000e-07 V_low
+ 6.386010000e-07 V_low
+ 6.387000000e-07 V_low
+ 6.387010000e-07 V_low
+ 6.388000000e-07 V_low
+ 6.388010000e-07 V_low
+ 6.389000000e-07 V_low
+ 6.389010000e-07 V_hig
+ 6.390000000e-07 V_hig
+ 6.390010000e-07 V_hig
+ 6.391000000e-07 V_hig
+ 6.391010000e-07 V_hig
+ 6.392000000e-07 V_hig
+ 6.392010000e-07 V_hig
+ 6.393000000e-07 V_hig
+ 6.393010000e-07 V_hig
+ 6.394000000e-07 V_hig
+ 6.394010000e-07 V_hig
+ 6.395000000e-07 V_hig
+ 6.395010000e-07 V_hig
+ 6.396000000e-07 V_hig
+ 6.396010000e-07 V_hig
+ 6.397000000e-07 V_hig
+ 6.397010000e-07 V_hig
+ 6.398000000e-07 V_hig
+ 6.398010000e-07 V_hig
+ 6.399000000e-07 V_hig
+ 6.399010000e-07 V_hig
+ 6.400000000e-07 V_hig
+ 6.400010000e-07 V_hig
+ 6.401000000e-07 V_hig
+ 6.401010000e-07 V_hig
+ 6.402000000e-07 V_hig
+ 6.402010000e-07 V_hig
+ 6.403000000e-07 V_hig
+ 6.403010000e-07 V_hig
+ 6.404000000e-07 V_hig
+ 6.404010000e-07 V_hig
+ 6.405000000e-07 V_hig
+ 6.405010000e-07 V_hig
+ 6.406000000e-07 V_hig
+ 6.406010000e-07 V_hig
+ 6.407000000e-07 V_hig
+ 6.407010000e-07 V_hig
+ 6.408000000e-07 V_hig
+ 6.408010000e-07 V_hig
+ 6.409000000e-07 V_hig
+ 6.409010000e-07 V_low
+ 6.410000000e-07 V_low
+ 6.410010000e-07 V_low
+ 6.411000000e-07 V_low
+ 6.411010000e-07 V_low
+ 6.412000000e-07 V_low
+ 6.412010000e-07 V_low
+ 6.413000000e-07 V_low
+ 6.413010000e-07 V_low
+ 6.414000000e-07 V_low
+ 6.414010000e-07 V_low
+ 6.415000000e-07 V_low
+ 6.415010000e-07 V_low
+ 6.416000000e-07 V_low
+ 6.416010000e-07 V_low
+ 6.417000000e-07 V_low
+ 6.417010000e-07 V_low
+ 6.418000000e-07 V_low
+ 6.418010000e-07 V_low
+ 6.419000000e-07 V_low
+ 6.419010000e-07 V_low
+ 6.420000000e-07 V_low
+ 6.420010000e-07 V_low
+ 6.421000000e-07 V_low
+ 6.421010000e-07 V_low
+ 6.422000000e-07 V_low
+ 6.422010000e-07 V_low
+ 6.423000000e-07 V_low
+ 6.423010000e-07 V_low
+ 6.424000000e-07 V_low
+ 6.424010000e-07 V_low
+ 6.425000000e-07 V_low
+ 6.425010000e-07 V_low
+ 6.426000000e-07 V_low
+ 6.426010000e-07 V_low
+ 6.427000000e-07 V_low
+ 6.427010000e-07 V_low
+ 6.428000000e-07 V_low
+ 6.428010000e-07 V_low
+ 6.429000000e-07 V_low
+ 6.429010000e-07 V_hig
+ 6.430000000e-07 V_hig
+ 6.430010000e-07 V_hig
+ 6.431000000e-07 V_hig
+ 6.431010000e-07 V_hig
+ 6.432000000e-07 V_hig
+ 6.432010000e-07 V_hig
+ 6.433000000e-07 V_hig
+ 6.433010000e-07 V_hig
+ 6.434000000e-07 V_hig
+ 6.434010000e-07 V_hig
+ 6.435000000e-07 V_hig
+ 6.435010000e-07 V_hig
+ 6.436000000e-07 V_hig
+ 6.436010000e-07 V_hig
+ 6.437000000e-07 V_hig
+ 6.437010000e-07 V_hig
+ 6.438000000e-07 V_hig
+ 6.438010000e-07 V_hig
+ 6.439000000e-07 V_hig
+ 6.439010000e-07 V_low
+ 6.440000000e-07 V_low
+ 6.440010000e-07 V_low
+ 6.441000000e-07 V_low
+ 6.441010000e-07 V_low
+ 6.442000000e-07 V_low
+ 6.442010000e-07 V_low
+ 6.443000000e-07 V_low
+ 6.443010000e-07 V_low
+ 6.444000000e-07 V_low
+ 6.444010000e-07 V_low
+ 6.445000000e-07 V_low
+ 6.445010000e-07 V_low
+ 6.446000000e-07 V_low
+ 6.446010000e-07 V_low
+ 6.447000000e-07 V_low
+ 6.447010000e-07 V_low
+ 6.448000000e-07 V_low
+ 6.448010000e-07 V_low
+ 6.449000000e-07 V_low
+ 6.449010000e-07 V_hig
+ 6.450000000e-07 V_hig
+ 6.450010000e-07 V_hig
+ 6.451000000e-07 V_hig
+ 6.451010000e-07 V_hig
+ 6.452000000e-07 V_hig
+ 6.452010000e-07 V_hig
+ 6.453000000e-07 V_hig
+ 6.453010000e-07 V_hig
+ 6.454000000e-07 V_hig
+ 6.454010000e-07 V_hig
+ 6.455000000e-07 V_hig
+ 6.455010000e-07 V_hig
+ 6.456000000e-07 V_hig
+ 6.456010000e-07 V_hig
+ 6.457000000e-07 V_hig
+ 6.457010000e-07 V_hig
+ 6.458000000e-07 V_hig
+ 6.458010000e-07 V_hig
+ 6.459000000e-07 V_hig
+ 6.459010000e-07 V_hig
+ 6.460000000e-07 V_hig
+ 6.460010000e-07 V_hig
+ 6.461000000e-07 V_hig
+ 6.461010000e-07 V_hig
+ 6.462000000e-07 V_hig
+ 6.462010000e-07 V_hig
+ 6.463000000e-07 V_hig
+ 6.463010000e-07 V_hig
+ 6.464000000e-07 V_hig
+ 6.464010000e-07 V_hig
+ 6.465000000e-07 V_hig
+ 6.465010000e-07 V_hig
+ 6.466000000e-07 V_hig
+ 6.466010000e-07 V_hig
+ 6.467000000e-07 V_hig
+ 6.467010000e-07 V_hig
+ 6.468000000e-07 V_hig
+ 6.468010000e-07 V_hig
+ 6.469000000e-07 V_hig
+ 6.469010000e-07 V_hig
+ 6.470000000e-07 V_hig
+ 6.470010000e-07 V_hig
+ 6.471000000e-07 V_hig
+ 6.471010000e-07 V_hig
+ 6.472000000e-07 V_hig
+ 6.472010000e-07 V_hig
+ 6.473000000e-07 V_hig
+ 6.473010000e-07 V_hig
+ 6.474000000e-07 V_hig
+ 6.474010000e-07 V_hig
+ 6.475000000e-07 V_hig
+ 6.475010000e-07 V_hig
+ 6.476000000e-07 V_hig
+ 6.476010000e-07 V_hig
+ 6.477000000e-07 V_hig
+ 6.477010000e-07 V_hig
+ 6.478000000e-07 V_hig
+ 6.478010000e-07 V_hig
+ 6.479000000e-07 V_hig
+ 6.479010000e-07 V_low
+ 6.480000000e-07 V_low
+ 6.480010000e-07 V_low
+ 6.481000000e-07 V_low
+ 6.481010000e-07 V_low
+ 6.482000000e-07 V_low
+ 6.482010000e-07 V_low
+ 6.483000000e-07 V_low
+ 6.483010000e-07 V_low
+ 6.484000000e-07 V_low
+ 6.484010000e-07 V_low
+ 6.485000000e-07 V_low
+ 6.485010000e-07 V_low
+ 6.486000000e-07 V_low
+ 6.486010000e-07 V_low
+ 6.487000000e-07 V_low
+ 6.487010000e-07 V_low
+ 6.488000000e-07 V_low
+ 6.488010000e-07 V_low
+ 6.489000000e-07 V_low
+ 6.489010000e-07 V_low
+ 6.490000000e-07 V_low
+ 6.490010000e-07 V_low
+ 6.491000000e-07 V_low
+ 6.491010000e-07 V_low
+ 6.492000000e-07 V_low
+ 6.492010000e-07 V_low
+ 6.493000000e-07 V_low
+ 6.493010000e-07 V_low
+ 6.494000000e-07 V_low
+ 6.494010000e-07 V_low
+ 6.495000000e-07 V_low
+ 6.495010000e-07 V_low
+ 6.496000000e-07 V_low
+ 6.496010000e-07 V_low
+ 6.497000000e-07 V_low
+ 6.497010000e-07 V_low
+ 6.498000000e-07 V_low
+ 6.498010000e-07 V_low
+ 6.499000000e-07 V_low
+ 6.499010000e-07 V_low
+ 6.500000000e-07 V_low
+ 6.500010000e-07 V_low
+ 6.501000000e-07 V_low
+ 6.501010000e-07 V_low
+ 6.502000000e-07 V_low
+ 6.502010000e-07 V_low
+ 6.503000000e-07 V_low
+ 6.503010000e-07 V_low
+ 6.504000000e-07 V_low
+ 6.504010000e-07 V_low
+ 6.505000000e-07 V_low
+ 6.505010000e-07 V_low
+ 6.506000000e-07 V_low
+ 6.506010000e-07 V_low
+ 6.507000000e-07 V_low
+ 6.507010000e-07 V_low
+ 6.508000000e-07 V_low
+ 6.508010000e-07 V_low
+ 6.509000000e-07 V_low
+ 6.509010000e-07 V_hig
+ 6.510000000e-07 V_hig
+ 6.510010000e-07 V_hig
+ 6.511000000e-07 V_hig
+ 6.511010000e-07 V_hig
+ 6.512000000e-07 V_hig
+ 6.512010000e-07 V_hig
+ 6.513000000e-07 V_hig
+ 6.513010000e-07 V_hig
+ 6.514000000e-07 V_hig
+ 6.514010000e-07 V_hig
+ 6.515000000e-07 V_hig
+ 6.515010000e-07 V_hig
+ 6.516000000e-07 V_hig
+ 6.516010000e-07 V_hig
+ 6.517000000e-07 V_hig
+ 6.517010000e-07 V_hig
+ 6.518000000e-07 V_hig
+ 6.518010000e-07 V_hig
+ 6.519000000e-07 V_hig
+ 6.519010000e-07 V_low
+ 6.520000000e-07 V_low
+ 6.520010000e-07 V_low
+ 6.521000000e-07 V_low
+ 6.521010000e-07 V_low
+ 6.522000000e-07 V_low
+ 6.522010000e-07 V_low
+ 6.523000000e-07 V_low
+ 6.523010000e-07 V_low
+ 6.524000000e-07 V_low
+ 6.524010000e-07 V_low
+ 6.525000000e-07 V_low
+ 6.525010000e-07 V_low
+ 6.526000000e-07 V_low
+ 6.526010000e-07 V_low
+ 6.527000000e-07 V_low
+ 6.527010000e-07 V_low
+ 6.528000000e-07 V_low
+ 6.528010000e-07 V_low
+ 6.529000000e-07 V_low
+ 6.529010000e-07 V_low
+ 6.530000000e-07 V_low
+ 6.530010000e-07 V_low
+ 6.531000000e-07 V_low
+ 6.531010000e-07 V_low
+ 6.532000000e-07 V_low
+ 6.532010000e-07 V_low
+ 6.533000000e-07 V_low
+ 6.533010000e-07 V_low
+ 6.534000000e-07 V_low
+ 6.534010000e-07 V_low
+ 6.535000000e-07 V_low
+ 6.535010000e-07 V_low
+ 6.536000000e-07 V_low
+ 6.536010000e-07 V_low
+ 6.537000000e-07 V_low
+ 6.537010000e-07 V_low
+ 6.538000000e-07 V_low
+ 6.538010000e-07 V_low
+ 6.539000000e-07 V_low
+ 6.539010000e-07 V_low
+ 6.540000000e-07 V_low
+ 6.540010000e-07 V_low
+ 6.541000000e-07 V_low
+ 6.541010000e-07 V_low
+ 6.542000000e-07 V_low
+ 6.542010000e-07 V_low
+ 6.543000000e-07 V_low
+ 6.543010000e-07 V_low
+ 6.544000000e-07 V_low
+ 6.544010000e-07 V_low
+ 6.545000000e-07 V_low
+ 6.545010000e-07 V_low
+ 6.546000000e-07 V_low
+ 6.546010000e-07 V_low
+ 6.547000000e-07 V_low
+ 6.547010000e-07 V_low
+ 6.548000000e-07 V_low
+ 6.548010000e-07 V_low
+ 6.549000000e-07 V_low
+ 6.549010000e-07 V_low
+ 6.550000000e-07 V_low
+ 6.550010000e-07 V_low
+ 6.551000000e-07 V_low
+ 6.551010000e-07 V_low
+ 6.552000000e-07 V_low
+ 6.552010000e-07 V_low
+ 6.553000000e-07 V_low
+ 6.553010000e-07 V_low
+ 6.554000000e-07 V_low
+ 6.554010000e-07 V_low
+ 6.555000000e-07 V_low
+ 6.555010000e-07 V_low
+ 6.556000000e-07 V_low
+ 6.556010000e-07 V_low
+ 6.557000000e-07 V_low
+ 6.557010000e-07 V_low
+ 6.558000000e-07 V_low
+ 6.558010000e-07 V_low
+ 6.559000000e-07 V_low
+ 6.559010000e-07 V_hig
+ 6.560000000e-07 V_hig
+ 6.560010000e-07 V_hig
+ 6.561000000e-07 V_hig
+ 6.561010000e-07 V_hig
+ 6.562000000e-07 V_hig
+ 6.562010000e-07 V_hig
+ 6.563000000e-07 V_hig
+ 6.563010000e-07 V_hig
+ 6.564000000e-07 V_hig
+ 6.564010000e-07 V_hig
+ 6.565000000e-07 V_hig
+ 6.565010000e-07 V_hig
+ 6.566000000e-07 V_hig
+ 6.566010000e-07 V_hig
+ 6.567000000e-07 V_hig
+ 6.567010000e-07 V_hig
+ 6.568000000e-07 V_hig
+ 6.568010000e-07 V_hig
+ 6.569000000e-07 V_hig
+ 6.569010000e-07 V_hig
+ 6.570000000e-07 V_hig
+ 6.570010000e-07 V_hig
+ 6.571000000e-07 V_hig
+ 6.571010000e-07 V_hig
+ 6.572000000e-07 V_hig
+ 6.572010000e-07 V_hig
+ 6.573000000e-07 V_hig
+ 6.573010000e-07 V_hig
+ 6.574000000e-07 V_hig
+ 6.574010000e-07 V_hig
+ 6.575000000e-07 V_hig
+ 6.575010000e-07 V_hig
+ 6.576000000e-07 V_hig
+ 6.576010000e-07 V_hig
+ 6.577000000e-07 V_hig
+ 6.577010000e-07 V_hig
+ 6.578000000e-07 V_hig
+ 6.578010000e-07 V_hig
+ 6.579000000e-07 V_hig
+ 6.579010000e-07 V_low
+ 6.580000000e-07 V_low
+ 6.580010000e-07 V_low
+ 6.581000000e-07 V_low
+ 6.581010000e-07 V_low
+ 6.582000000e-07 V_low
+ 6.582010000e-07 V_low
+ 6.583000000e-07 V_low
+ 6.583010000e-07 V_low
+ 6.584000000e-07 V_low
+ 6.584010000e-07 V_low
+ 6.585000000e-07 V_low
+ 6.585010000e-07 V_low
+ 6.586000000e-07 V_low
+ 6.586010000e-07 V_low
+ 6.587000000e-07 V_low
+ 6.587010000e-07 V_low
+ 6.588000000e-07 V_low
+ 6.588010000e-07 V_low
+ 6.589000000e-07 V_low
+ 6.589010000e-07 V_low
+ 6.590000000e-07 V_low
+ 6.590010000e-07 V_low
+ 6.591000000e-07 V_low
+ 6.591010000e-07 V_low
+ 6.592000000e-07 V_low
+ 6.592010000e-07 V_low
+ 6.593000000e-07 V_low
+ 6.593010000e-07 V_low
+ 6.594000000e-07 V_low
+ 6.594010000e-07 V_low
+ 6.595000000e-07 V_low
+ 6.595010000e-07 V_low
+ 6.596000000e-07 V_low
+ 6.596010000e-07 V_low
+ 6.597000000e-07 V_low
+ 6.597010000e-07 V_low
+ 6.598000000e-07 V_low
+ 6.598010000e-07 V_low
+ 6.599000000e-07 V_low
+ 6.599010000e-07 V_hig
+ 6.600000000e-07 V_hig
+ 6.600010000e-07 V_hig
+ 6.601000000e-07 V_hig
+ 6.601010000e-07 V_hig
+ 6.602000000e-07 V_hig
+ 6.602010000e-07 V_hig
+ 6.603000000e-07 V_hig
+ 6.603010000e-07 V_hig
+ 6.604000000e-07 V_hig
+ 6.604010000e-07 V_hig
+ 6.605000000e-07 V_hig
+ 6.605010000e-07 V_hig
+ 6.606000000e-07 V_hig
+ 6.606010000e-07 V_hig
+ 6.607000000e-07 V_hig
+ 6.607010000e-07 V_hig
+ 6.608000000e-07 V_hig
+ 6.608010000e-07 V_hig
+ 6.609000000e-07 V_hig
+ 6.609010000e-07 V_low
+ 6.610000000e-07 V_low
+ 6.610010000e-07 V_low
+ 6.611000000e-07 V_low
+ 6.611010000e-07 V_low
+ 6.612000000e-07 V_low
+ 6.612010000e-07 V_low
+ 6.613000000e-07 V_low
+ 6.613010000e-07 V_low
+ 6.614000000e-07 V_low
+ 6.614010000e-07 V_low
+ 6.615000000e-07 V_low
+ 6.615010000e-07 V_low
+ 6.616000000e-07 V_low
+ 6.616010000e-07 V_low
+ 6.617000000e-07 V_low
+ 6.617010000e-07 V_low
+ 6.618000000e-07 V_low
+ 6.618010000e-07 V_low
+ 6.619000000e-07 V_low
+ 6.619010000e-07 V_low
+ 6.620000000e-07 V_low
+ 6.620010000e-07 V_low
+ 6.621000000e-07 V_low
+ 6.621010000e-07 V_low
+ 6.622000000e-07 V_low
+ 6.622010000e-07 V_low
+ 6.623000000e-07 V_low
+ 6.623010000e-07 V_low
+ 6.624000000e-07 V_low
+ 6.624010000e-07 V_low
+ 6.625000000e-07 V_low
+ 6.625010000e-07 V_low
+ 6.626000000e-07 V_low
+ 6.626010000e-07 V_low
+ 6.627000000e-07 V_low
+ 6.627010000e-07 V_low
+ 6.628000000e-07 V_low
+ 6.628010000e-07 V_low
+ 6.629000000e-07 V_low
+ 6.629010000e-07 V_low
+ 6.630000000e-07 V_low
+ 6.630010000e-07 V_low
+ 6.631000000e-07 V_low
+ 6.631010000e-07 V_low
+ 6.632000000e-07 V_low
+ 6.632010000e-07 V_low
+ 6.633000000e-07 V_low
+ 6.633010000e-07 V_low
+ 6.634000000e-07 V_low
+ 6.634010000e-07 V_low
+ 6.635000000e-07 V_low
+ 6.635010000e-07 V_low
+ 6.636000000e-07 V_low
+ 6.636010000e-07 V_low
+ 6.637000000e-07 V_low
+ 6.637010000e-07 V_low
+ 6.638000000e-07 V_low
+ 6.638010000e-07 V_low
+ 6.639000000e-07 V_low
+ 6.639010000e-07 V_hig
+ 6.640000000e-07 V_hig
+ 6.640010000e-07 V_hig
+ 6.641000000e-07 V_hig
+ 6.641010000e-07 V_hig
+ 6.642000000e-07 V_hig
+ 6.642010000e-07 V_hig
+ 6.643000000e-07 V_hig
+ 6.643010000e-07 V_hig
+ 6.644000000e-07 V_hig
+ 6.644010000e-07 V_hig
+ 6.645000000e-07 V_hig
+ 6.645010000e-07 V_hig
+ 6.646000000e-07 V_hig
+ 6.646010000e-07 V_hig
+ 6.647000000e-07 V_hig
+ 6.647010000e-07 V_hig
+ 6.648000000e-07 V_hig
+ 6.648010000e-07 V_hig
+ 6.649000000e-07 V_hig
+ 6.649010000e-07 V_low
+ 6.650000000e-07 V_low
+ 6.650010000e-07 V_low
+ 6.651000000e-07 V_low
+ 6.651010000e-07 V_low
+ 6.652000000e-07 V_low
+ 6.652010000e-07 V_low
+ 6.653000000e-07 V_low
+ 6.653010000e-07 V_low
+ 6.654000000e-07 V_low
+ 6.654010000e-07 V_low
+ 6.655000000e-07 V_low
+ 6.655010000e-07 V_low
+ 6.656000000e-07 V_low
+ 6.656010000e-07 V_low
+ 6.657000000e-07 V_low
+ 6.657010000e-07 V_low
+ 6.658000000e-07 V_low
+ 6.658010000e-07 V_low
+ 6.659000000e-07 V_low
+ 6.659010000e-07 V_hig
+ 6.660000000e-07 V_hig
+ 6.660010000e-07 V_hig
+ 6.661000000e-07 V_hig
+ 6.661010000e-07 V_hig
+ 6.662000000e-07 V_hig
+ 6.662010000e-07 V_hig
+ 6.663000000e-07 V_hig
+ 6.663010000e-07 V_hig
+ 6.664000000e-07 V_hig
+ 6.664010000e-07 V_hig
+ 6.665000000e-07 V_hig
+ 6.665010000e-07 V_hig
+ 6.666000000e-07 V_hig
+ 6.666010000e-07 V_hig
+ 6.667000000e-07 V_hig
+ 6.667010000e-07 V_hig
+ 6.668000000e-07 V_hig
+ 6.668010000e-07 V_hig
+ 6.669000000e-07 V_hig
+ 6.669010000e-07 V_low
+ 6.670000000e-07 V_low
+ 6.670010000e-07 V_low
+ 6.671000000e-07 V_low
+ 6.671010000e-07 V_low
+ 6.672000000e-07 V_low
+ 6.672010000e-07 V_low
+ 6.673000000e-07 V_low
+ 6.673010000e-07 V_low
+ 6.674000000e-07 V_low
+ 6.674010000e-07 V_low
+ 6.675000000e-07 V_low
+ 6.675010000e-07 V_low
+ 6.676000000e-07 V_low
+ 6.676010000e-07 V_low
+ 6.677000000e-07 V_low
+ 6.677010000e-07 V_low
+ 6.678000000e-07 V_low
+ 6.678010000e-07 V_low
+ 6.679000000e-07 V_low
+ 6.679010000e-07 V_low
+ 6.680000000e-07 V_low
+ 6.680010000e-07 V_low
+ 6.681000000e-07 V_low
+ 6.681010000e-07 V_low
+ 6.682000000e-07 V_low
+ 6.682010000e-07 V_low
+ 6.683000000e-07 V_low
+ 6.683010000e-07 V_low
+ 6.684000000e-07 V_low
+ 6.684010000e-07 V_low
+ 6.685000000e-07 V_low
+ 6.685010000e-07 V_low
+ 6.686000000e-07 V_low
+ 6.686010000e-07 V_low
+ 6.687000000e-07 V_low
+ 6.687010000e-07 V_low
+ 6.688000000e-07 V_low
+ 6.688010000e-07 V_low
+ 6.689000000e-07 V_low
+ 6.689010000e-07 V_hig
+ 6.690000000e-07 V_hig
+ 6.690010000e-07 V_hig
+ 6.691000000e-07 V_hig
+ 6.691010000e-07 V_hig
+ 6.692000000e-07 V_hig
+ 6.692010000e-07 V_hig
+ 6.693000000e-07 V_hig
+ 6.693010000e-07 V_hig
+ 6.694000000e-07 V_hig
+ 6.694010000e-07 V_hig
+ 6.695000000e-07 V_hig
+ 6.695010000e-07 V_hig
+ 6.696000000e-07 V_hig
+ 6.696010000e-07 V_hig
+ 6.697000000e-07 V_hig
+ 6.697010000e-07 V_hig
+ 6.698000000e-07 V_hig
+ 6.698010000e-07 V_hig
+ 6.699000000e-07 V_hig
+ 6.699010000e-07 V_low
+ 6.700000000e-07 V_low
+ 6.700010000e-07 V_low
+ 6.701000000e-07 V_low
+ 6.701010000e-07 V_low
+ 6.702000000e-07 V_low
+ 6.702010000e-07 V_low
+ 6.703000000e-07 V_low
+ 6.703010000e-07 V_low
+ 6.704000000e-07 V_low
+ 6.704010000e-07 V_low
+ 6.705000000e-07 V_low
+ 6.705010000e-07 V_low
+ 6.706000000e-07 V_low
+ 6.706010000e-07 V_low
+ 6.707000000e-07 V_low
+ 6.707010000e-07 V_low
+ 6.708000000e-07 V_low
+ 6.708010000e-07 V_low
+ 6.709000000e-07 V_low
+ 6.709010000e-07 V_low
+ 6.710000000e-07 V_low
+ 6.710010000e-07 V_low
+ 6.711000000e-07 V_low
+ 6.711010000e-07 V_low
+ 6.712000000e-07 V_low
+ 6.712010000e-07 V_low
+ 6.713000000e-07 V_low
+ 6.713010000e-07 V_low
+ 6.714000000e-07 V_low
+ 6.714010000e-07 V_low
+ 6.715000000e-07 V_low
+ 6.715010000e-07 V_low
+ 6.716000000e-07 V_low
+ 6.716010000e-07 V_low
+ 6.717000000e-07 V_low
+ 6.717010000e-07 V_low
+ 6.718000000e-07 V_low
+ 6.718010000e-07 V_low
+ 6.719000000e-07 V_low
+ 6.719010000e-07 V_hig
+ 6.720000000e-07 V_hig
+ 6.720010000e-07 V_hig
+ 6.721000000e-07 V_hig
+ 6.721010000e-07 V_hig
+ 6.722000000e-07 V_hig
+ 6.722010000e-07 V_hig
+ 6.723000000e-07 V_hig
+ 6.723010000e-07 V_hig
+ 6.724000000e-07 V_hig
+ 6.724010000e-07 V_hig
+ 6.725000000e-07 V_hig
+ 6.725010000e-07 V_hig
+ 6.726000000e-07 V_hig
+ 6.726010000e-07 V_hig
+ 6.727000000e-07 V_hig
+ 6.727010000e-07 V_hig
+ 6.728000000e-07 V_hig
+ 6.728010000e-07 V_hig
+ 6.729000000e-07 V_hig
+ 6.729010000e-07 V_hig
+ 6.730000000e-07 V_hig
+ 6.730010000e-07 V_hig
+ 6.731000000e-07 V_hig
+ 6.731010000e-07 V_hig
+ 6.732000000e-07 V_hig
+ 6.732010000e-07 V_hig
+ 6.733000000e-07 V_hig
+ 6.733010000e-07 V_hig
+ 6.734000000e-07 V_hig
+ 6.734010000e-07 V_hig
+ 6.735000000e-07 V_hig
+ 6.735010000e-07 V_hig
+ 6.736000000e-07 V_hig
+ 6.736010000e-07 V_hig
+ 6.737000000e-07 V_hig
+ 6.737010000e-07 V_hig
+ 6.738000000e-07 V_hig
+ 6.738010000e-07 V_hig
+ 6.739000000e-07 V_hig
+ 6.739010000e-07 V_low
+ 6.740000000e-07 V_low
+ 6.740010000e-07 V_low
+ 6.741000000e-07 V_low
+ 6.741010000e-07 V_low
+ 6.742000000e-07 V_low
+ 6.742010000e-07 V_low
+ 6.743000000e-07 V_low
+ 6.743010000e-07 V_low
+ 6.744000000e-07 V_low
+ 6.744010000e-07 V_low
+ 6.745000000e-07 V_low
+ 6.745010000e-07 V_low
+ 6.746000000e-07 V_low
+ 6.746010000e-07 V_low
+ 6.747000000e-07 V_low
+ 6.747010000e-07 V_low
+ 6.748000000e-07 V_low
+ 6.748010000e-07 V_low
+ 6.749000000e-07 V_low
+ 6.749010000e-07 V_low
+ 6.750000000e-07 V_low
+ 6.750010000e-07 V_low
+ 6.751000000e-07 V_low
+ 6.751010000e-07 V_low
+ 6.752000000e-07 V_low
+ 6.752010000e-07 V_low
+ 6.753000000e-07 V_low
+ 6.753010000e-07 V_low
+ 6.754000000e-07 V_low
+ 6.754010000e-07 V_low
+ 6.755000000e-07 V_low
+ 6.755010000e-07 V_low
+ 6.756000000e-07 V_low
+ 6.756010000e-07 V_low
+ 6.757000000e-07 V_low
+ 6.757010000e-07 V_low
+ 6.758000000e-07 V_low
+ 6.758010000e-07 V_low
+ 6.759000000e-07 V_low
+ 6.759010000e-07 V_low
+ 6.760000000e-07 V_low
+ 6.760010000e-07 V_low
+ 6.761000000e-07 V_low
+ 6.761010000e-07 V_low
+ 6.762000000e-07 V_low
+ 6.762010000e-07 V_low
+ 6.763000000e-07 V_low
+ 6.763010000e-07 V_low
+ 6.764000000e-07 V_low
+ 6.764010000e-07 V_low
+ 6.765000000e-07 V_low
+ 6.765010000e-07 V_low
+ 6.766000000e-07 V_low
+ 6.766010000e-07 V_low
+ 6.767000000e-07 V_low
+ 6.767010000e-07 V_low
+ 6.768000000e-07 V_low
+ 6.768010000e-07 V_low
+ 6.769000000e-07 V_low
+ 6.769010000e-07 V_low
+ 6.770000000e-07 V_low
+ 6.770010000e-07 V_low
+ 6.771000000e-07 V_low
+ 6.771010000e-07 V_low
+ 6.772000000e-07 V_low
+ 6.772010000e-07 V_low
+ 6.773000000e-07 V_low
+ 6.773010000e-07 V_low
+ 6.774000000e-07 V_low
+ 6.774010000e-07 V_low
+ 6.775000000e-07 V_low
+ 6.775010000e-07 V_low
+ 6.776000000e-07 V_low
+ 6.776010000e-07 V_low
+ 6.777000000e-07 V_low
+ 6.777010000e-07 V_low
+ 6.778000000e-07 V_low
+ 6.778010000e-07 V_low
+ 6.779000000e-07 V_low
+ 6.779010000e-07 V_hig
+ 6.780000000e-07 V_hig
+ 6.780010000e-07 V_hig
+ 6.781000000e-07 V_hig
+ 6.781010000e-07 V_hig
+ 6.782000000e-07 V_hig
+ 6.782010000e-07 V_hig
+ 6.783000000e-07 V_hig
+ 6.783010000e-07 V_hig
+ 6.784000000e-07 V_hig
+ 6.784010000e-07 V_hig
+ 6.785000000e-07 V_hig
+ 6.785010000e-07 V_hig
+ 6.786000000e-07 V_hig
+ 6.786010000e-07 V_hig
+ 6.787000000e-07 V_hig
+ 6.787010000e-07 V_hig
+ 6.788000000e-07 V_hig
+ 6.788010000e-07 V_hig
+ 6.789000000e-07 V_hig
+ 6.789010000e-07 V_hig
+ 6.790000000e-07 V_hig
+ 6.790010000e-07 V_hig
+ 6.791000000e-07 V_hig
+ 6.791010000e-07 V_hig
+ 6.792000000e-07 V_hig
+ 6.792010000e-07 V_hig
+ 6.793000000e-07 V_hig
+ 6.793010000e-07 V_hig
+ 6.794000000e-07 V_hig
+ 6.794010000e-07 V_hig
+ 6.795000000e-07 V_hig
+ 6.795010000e-07 V_hig
+ 6.796000000e-07 V_hig
+ 6.796010000e-07 V_hig
+ 6.797000000e-07 V_hig
+ 6.797010000e-07 V_hig
+ 6.798000000e-07 V_hig
+ 6.798010000e-07 V_hig
+ 6.799000000e-07 V_hig
+ 6.799010000e-07 V_hig
+ 6.800000000e-07 V_hig
+ 6.800010000e-07 V_hig
+ 6.801000000e-07 V_hig
+ 6.801010000e-07 V_hig
+ 6.802000000e-07 V_hig
+ 6.802010000e-07 V_hig
+ 6.803000000e-07 V_hig
+ 6.803010000e-07 V_hig
+ 6.804000000e-07 V_hig
+ 6.804010000e-07 V_hig
+ 6.805000000e-07 V_hig
+ 6.805010000e-07 V_hig
+ 6.806000000e-07 V_hig
+ 6.806010000e-07 V_hig
+ 6.807000000e-07 V_hig
+ 6.807010000e-07 V_hig
+ 6.808000000e-07 V_hig
+ 6.808010000e-07 V_hig
+ 6.809000000e-07 V_hig
+ 6.809010000e-07 V_hig
+ 6.810000000e-07 V_hig
+ 6.810010000e-07 V_hig
+ 6.811000000e-07 V_hig
+ 6.811010000e-07 V_hig
+ 6.812000000e-07 V_hig
+ 6.812010000e-07 V_hig
+ 6.813000000e-07 V_hig
+ 6.813010000e-07 V_hig
+ 6.814000000e-07 V_hig
+ 6.814010000e-07 V_hig
+ 6.815000000e-07 V_hig
+ 6.815010000e-07 V_hig
+ 6.816000000e-07 V_hig
+ 6.816010000e-07 V_hig
+ 6.817000000e-07 V_hig
+ 6.817010000e-07 V_hig
+ 6.818000000e-07 V_hig
+ 6.818010000e-07 V_hig
+ 6.819000000e-07 V_hig
+ 6.819010000e-07 V_low
+ 6.820000000e-07 V_low
+ 6.820010000e-07 V_low
+ 6.821000000e-07 V_low
+ 6.821010000e-07 V_low
+ 6.822000000e-07 V_low
+ 6.822010000e-07 V_low
+ 6.823000000e-07 V_low
+ 6.823010000e-07 V_low
+ 6.824000000e-07 V_low
+ 6.824010000e-07 V_low
+ 6.825000000e-07 V_low
+ 6.825010000e-07 V_low
+ 6.826000000e-07 V_low
+ 6.826010000e-07 V_low
+ 6.827000000e-07 V_low
+ 6.827010000e-07 V_low
+ 6.828000000e-07 V_low
+ 6.828010000e-07 V_low
+ 6.829000000e-07 V_low
+ 6.829010000e-07 V_hig
+ 6.830000000e-07 V_hig
+ 6.830010000e-07 V_hig
+ 6.831000000e-07 V_hig
+ 6.831010000e-07 V_hig
+ 6.832000000e-07 V_hig
+ 6.832010000e-07 V_hig
+ 6.833000000e-07 V_hig
+ 6.833010000e-07 V_hig
+ 6.834000000e-07 V_hig
+ 6.834010000e-07 V_hig
+ 6.835000000e-07 V_hig
+ 6.835010000e-07 V_hig
+ 6.836000000e-07 V_hig
+ 6.836010000e-07 V_hig
+ 6.837000000e-07 V_hig
+ 6.837010000e-07 V_hig
+ 6.838000000e-07 V_hig
+ 6.838010000e-07 V_hig
+ 6.839000000e-07 V_hig
+ 6.839010000e-07 V_hig
+ 6.840000000e-07 V_hig
+ 6.840010000e-07 V_hig
+ 6.841000000e-07 V_hig
+ 6.841010000e-07 V_hig
+ 6.842000000e-07 V_hig
+ 6.842010000e-07 V_hig
+ 6.843000000e-07 V_hig
+ 6.843010000e-07 V_hig
+ 6.844000000e-07 V_hig
+ 6.844010000e-07 V_hig
+ 6.845000000e-07 V_hig
+ 6.845010000e-07 V_hig
+ 6.846000000e-07 V_hig
+ 6.846010000e-07 V_hig
+ 6.847000000e-07 V_hig
+ 6.847010000e-07 V_hig
+ 6.848000000e-07 V_hig
+ 6.848010000e-07 V_hig
+ 6.849000000e-07 V_hig
+ 6.849010000e-07 V_low
+ 6.850000000e-07 V_low
+ 6.850010000e-07 V_low
+ 6.851000000e-07 V_low
+ 6.851010000e-07 V_low
+ 6.852000000e-07 V_low
+ 6.852010000e-07 V_low
+ 6.853000000e-07 V_low
+ 6.853010000e-07 V_low
+ 6.854000000e-07 V_low
+ 6.854010000e-07 V_low
+ 6.855000000e-07 V_low
+ 6.855010000e-07 V_low
+ 6.856000000e-07 V_low
+ 6.856010000e-07 V_low
+ 6.857000000e-07 V_low
+ 6.857010000e-07 V_low
+ 6.858000000e-07 V_low
+ 6.858010000e-07 V_low
+ 6.859000000e-07 V_low
+ 6.859010000e-07 V_low
+ 6.860000000e-07 V_low
+ 6.860010000e-07 V_low
+ 6.861000000e-07 V_low
+ 6.861010000e-07 V_low
+ 6.862000000e-07 V_low
+ 6.862010000e-07 V_low
+ 6.863000000e-07 V_low
+ 6.863010000e-07 V_low
+ 6.864000000e-07 V_low
+ 6.864010000e-07 V_low
+ 6.865000000e-07 V_low
+ 6.865010000e-07 V_low
+ 6.866000000e-07 V_low
+ 6.866010000e-07 V_low
+ 6.867000000e-07 V_low
+ 6.867010000e-07 V_low
+ 6.868000000e-07 V_low
+ 6.868010000e-07 V_low
+ 6.869000000e-07 V_low
+ 6.869010000e-07 V_hig
+ 6.870000000e-07 V_hig
+ 6.870010000e-07 V_hig
+ 6.871000000e-07 V_hig
+ 6.871010000e-07 V_hig
+ 6.872000000e-07 V_hig
+ 6.872010000e-07 V_hig
+ 6.873000000e-07 V_hig
+ 6.873010000e-07 V_hig
+ 6.874000000e-07 V_hig
+ 6.874010000e-07 V_hig
+ 6.875000000e-07 V_hig
+ 6.875010000e-07 V_hig
+ 6.876000000e-07 V_hig
+ 6.876010000e-07 V_hig
+ 6.877000000e-07 V_hig
+ 6.877010000e-07 V_hig
+ 6.878000000e-07 V_hig
+ 6.878010000e-07 V_hig
+ 6.879000000e-07 V_hig
+ 6.879010000e-07 V_hig
+ 6.880000000e-07 V_hig
+ 6.880010000e-07 V_hig
+ 6.881000000e-07 V_hig
+ 6.881010000e-07 V_hig
+ 6.882000000e-07 V_hig
+ 6.882010000e-07 V_hig
+ 6.883000000e-07 V_hig
+ 6.883010000e-07 V_hig
+ 6.884000000e-07 V_hig
+ 6.884010000e-07 V_hig
+ 6.885000000e-07 V_hig
+ 6.885010000e-07 V_hig
+ 6.886000000e-07 V_hig
+ 6.886010000e-07 V_hig
+ 6.887000000e-07 V_hig
+ 6.887010000e-07 V_hig
+ 6.888000000e-07 V_hig
+ 6.888010000e-07 V_hig
+ 6.889000000e-07 V_hig
+ 6.889010000e-07 V_low
+ 6.890000000e-07 V_low
+ 6.890010000e-07 V_low
+ 6.891000000e-07 V_low
+ 6.891010000e-07 V_low
+ 6.892000000e-07 V_low
+ 6.892010000e-07 V_low
+ 6.893000000e-07 V_low
+ 6.893010000e-07 V_low
+ 6.894000000e-07 V_low
+ 6.894010000e-07 V_low
+ 6.895000000e-07 V_low
+ 6.895010000e-07 V_low
+ 6.896000000e-07 V_low
+ 6.896010000e-07 V_low
+ 6.897000000e-07 V_low
+ 6.897010000e-07 V_low
+ 6.898000000e-07 V_low
+ 6.898010000e-07 V_low
+ 6.899000000e-07 V_low
+ 6.899010000e-07 V_hig
+ 6.900000000e-07 V_hig
+ 6.900010000e-07 V_hig
+ 6.901000000e-07 V_hig
+ 6.901010000e-07 V_hig
+ 6.902000000e-07 V_hig
+ 6.902010000e-07 V_hig
+ 6.903000000e-07 V_hig
+ 6.903010000e-07 V_hig
+ 6.904000000e-07 V_hig
+ 6.904010000e-07 V_hig
+ 6.905000000e-07 V_hig
+ 6.905010000e-07 V_hig
+ 6.906000000e-07 V_hig
+ 6.906010000e-07 V_hig
+ 6.907000000e-07 V_hig
+ 6.907010000e-07 V_hig
+ 6.908000000e-07 V_hig
+ 6.908010000e-07 V_hig
+ 6.909000000e-07 V_hig
+ 6.909010000e-07 V_hig
+ 6.910000000e-07 V_hig
+ 6.910010000e-07 V_hig
+ 6.911000000e-07 V_hig
+ 6.911010000e-07 V_hig
+ 6.912000000e-07 V_hig
+ 6.912010000e-07 V_hig
+ 6.913000000e-07 V_hig
+ 6.913010000e-07 V_hig
+ 6.914000000e-07 V_hig
+ 6.914010000e-07 V_hig
+ 6.915000000e-07 V_hig
+ 6.915010000e-07 V_hig
+ 6.916000000e-07 V_hig
+ 6.916010000e-07 V_hig
+ 6.917000000e-07 V_hig
+ 6.917010000e-07 V_hig
+ 6.918000000e-07 V_hig
+ 6.918010000e-07 V_hig
+ 6.919000000e-07 V_hig
+ 6.919010000e-07 V_low
+ 6.920000000e-07 V_low
+ 6.920010000e-07 V_low
+ 6.921000000e-07 V_low
+ 6.921010000e-07 V_low
+ 6.922000000e-07 V_low
+ 6.922010000e-07 V_low
+ 6.923000000e-07 V_low
+ 6.923010000e-07 V_low
+ 6.924000000e-07 V_low
+ 6.924010000e-07 V_low
+ 6.925000000e-07 V_low
+ 6.925010000e-07 V_low
+ 6.926000000e-07 V_low
+ 6.926010000e-07 V_low
+ 6.927000000e-07 V_low
+ 6.927010000e-07 V_low
+ 6.928000000e-07 V_low
+ 6.928010000e-07 V_low
+ 6.929000000e-07 V_low
+ 6.929010000e-07 V_low
+ 6.930000000e-07 V_low
+ 6.930010000e-07 V_low
+ 6.931000000e-07 V_low
+ 6.931010000e-07 V_low
+ 6.932000000e-07 V_low
+ 6.932010000e-07 V_low
+ 6.933000000e-07 V_low
+ 6.933010000e-07 V_low
+ 6.934000000e-07 V_low
+ 6.934010000e-07 V_low
+ 6.935000000e-07 V_low
+ 6.935010000e-07 V_low
+ 6.936000000e-07 V_low
+ 6.936010000e-07 V_low
+ 6.937000000e-07 V_low
+ 6.937010000e-07 V_low
+ 6.938000000e-07 V_low
+ 6.938010000e-07 V_low
+ 6.939000000e-07 V_low
+ 6.939010000e-07 V_low
+ 6.940000000e-07 V_low
+ 6.940010000e-07 V_low
+ 6.941000000e-07 V_low
+ 6.941010000e-07 V_low
+ 6.942000000e-07 V_low
+ 6.942010000e-07 V_low
+ 6.943000000e-07 V_low
+ 6.943010000e-07 V_low
+ 6.944000000e-07 V_low
+ 6.944010000e-07 V_low
+ 6.945000000e-07 V_low
+ 6.945010000e-07 V_low
+ 6.946000000e-07 V_low
+ 6.946010000e-07 V_low
+ 6.947000000e-07 V_low
+ 6.947010000e-07 V_low
+ 6.948000000e-07 V_low
+ 6.948010000e-07 V_low
+ 6.949000000e-07 V_low
+ 6.949010000e-07 V_low
+ 6.950000000e-07 V_low
+ 6.950010000e-07 V_low
+ 6.951000000e-07 V_low
+ 6.951010000e-07 V_low
+ 6.952000000e-07 V_low
+ 6.952010000e-07 V_low
+ 6.953000000e-07 V_low
+ 6.953010000e-07 V_low
+ 6.954000000e-07 V_low
+ 6.954010000e-07 V_low
+ 6.955000000e-07 V_low
+ 6.955010000e-07 V_low
+ 6.956000000e-07 V_low
+ 6.956010000e-07 V_low
+ 6.957000000e-07 V_low
+ 6.957010000e-07 V_low
+ 6.958000000e-07 V_low
+ 6.958010000e-07 V_low
+ 6.959000000e-07 V_low
+ 6.959010000e-07 V_hig
+ 6.960000000e-07 V_hig
+ 6.960010000e-07 V_hig
+ 6.961000000e-07 V_hig
+ 6.961010000e-07 V_hig
+ 6.962000000e-07 V_hig
+ 6.962010000e-07 V_hig
+ 6.963000000e-07 V_hig
+ 6.963010000e-07 V_hig
+ 6.964000000e-07 V_hig
+ 6.964010000e-07 V_hig
+ 6.965000000e-07 V_hig
+ 6.965010000e-07 V_hig
+ 6.966000000e-07 V_hig
+ 6.966010000e-07 V_hig
+ 6.967000000e-07 V_hig
+ 6.967010000e-07 V_hig
+ 6.968000000e-07 V_hig
+ 6.968010000e-07 V_hig
+ 6.969000000e-07 V_hig
+ 6.969010000e-07 V_hig
+ 6.970000000e-07 V_hig
+ 6.970010000e-07 V_hig
+ 6.971000000e-07 V_hig
+ 6.971010000e-07 V_hig
+ 6.972000000e-07 V_hig
+ 6.972010000e-07 V_hig
+ 6.973000000e-07 V_hig
+ 6.973010000e-07 V_hig
+ 6.974000000e-07 V_hig
+ 6.974010000e-07 V_hig
+ 6.975000000e-07 V_hig
+ 6.975010000e-07 V_hig
+ 6.976000000e-07 V_hig
+ 6.976010000e-07 V_hig
+ 6.977000000e-07 V_hig
+ 6.977010000e-07 V_hig
+ 6.978000000e-07 V_hig
+ 6.978010000e-07 V_hig
+ 6.979000000e-07 V_hig
+ 6.979010000e-07 V_low
+ 6.980000000e-07 V_low
+ 6.980010000e-07 V_low
+ 6.981000000e-07 V_low
+ 6.981010000e-07 V_low
+ 6.982000000e-07 V_low
+ 6.982010000e-07 V_low
+ 6.983000000e-07 V_low
+ 6.983010000e-07 V_low
+ 6.984000000e-07 V_low
+ 6.984010000e-07 V_low
+ 6.985000000e-07 V_low
+ 6.985010000e-07 V_low
+ 6.986000000e-07 V_low
+ 6.986010000e-07 V_low
+ 6.987000000e-07 V_low
+ 6.987010000e-07 V_low
+ 6.988000000e-07 V_low
+ 6.988010000e-07 V_low
+ 6.989000000e-07 V_low
+ 6.989010000e-07 V_hig
+ 6.990000000e-07 V_hig
+ 6.990010000e-07 V_hig
+ 6.991000000e-07 V_hig
+ 6.991010000e-07 V_hig
+ 6.992000000e-07 V_hig
+ 6.992010000e-07 V_hig
+ 6.993000000e-07 V_hig
+ 6.993010000e-07 V_hig
+ 6.994000000e-07 V_hig
+ 6.994010000e-07 V_hig
+ 6.995000000e-07 V_hig
+ 6.995010000e-07 V_hig
+ 6.996000000e-07 V_hig
+ 6.996010000e-07 V_hig
+ 6.997000000e-07 V_hig
+ 6.997010000e-07 V_hig
+ 6.998000000e-07 V_hig
+ 6.998010000e-07 V_hig
+ 6.999000000e-07 V_hig
+ 6.999010000e-07 V_hig
+ 7.000000000e-07 V_hig
+ 7.000010000e-07 V_hig
+ 7.001000000e-07 V_hig
+ 7.001010000e-07 V_hig
+ 7.002000000e-07 V_hig
+ 7.002010000e-07 V_hig
+ 7.003000000e-07 V_hig
+ 7.003010000e-07 V_hig
+ 7.004000000e-07 V_hig
+ 7.004010000e-07 V_hig
+ 7.005000000e-07 V_hig
+ 7.005010000e-07 V_hig
+ 7.006000000e-07 V_hig
+ 7.006010000e-07 V_hig
+ 7.007000000e-07 V_hig
+ 7.007010000e-07 V_hig
+ 7.008000000e-07 V_hig
+ 7.008010000e-07 V_hig
+ 7.009000000e-07 V_hig
+ 7.009010000e-07 V_hig
+ 7.010000000e-07 V_hig
+ 7.010010000e-07 V_hig
+ 7.011000000e-07 V_hig
+ 7.011010000e-07 V_hig
+ 7.012000000e-07 V_hig
+ 7.012010000e-07 V_hig
+ 7.013000000e-07 V_hig
+ 7.013010000e-07 V_hig
+ 7.014000000e-07 V_hig
+ 7.014010000e-07 V_hig
+ 7.015000000e-07 V_hig
+ 7.015010000e-07 V_hig
+ 7.016000000e-07 V_hig
+ 7.016010000e-07 V_hig
+ 7.017000000e-07 V_hig
+ 7.017010000e-07 V_hig
+ 7.018000000e-07 V_hig
+ 7.018010000e-07 V_hig
+ 7.019000000e-07 V_hig
+ 7.019010000e-07 V_hig
+ 7.020000000e-07 V_hig
+ 7.020010000e-07 V_hig
+ 7.021000000e-07 V_hig
+ 7.021010000e-07 V_hig
+ 7.022000000e-07 V_hig
+ 7.022010000e-07 V_hig
+ 7.023000000e-07 V_hig
+ 7.023010000e-07 V_hig
+ 7.024000000e-07 V_hig
+ 7.024010000e-07 V_hig
+ 7.025000000e-07 V_hig
+ 7.025010000e-07 V_hig
+ 7.026000000e-07 V_hig
+ 7.026010000e-07 V_hig
+ 7.027000000e-07 V_hig
+ 7.027010000e-07 V_hig
+ 7.028000000e-07 V_hig
+ 7.028010000e-07 V_hig
+ 7.029000000e-07 V_hig
+ 7.029010000e-07 V_low
+ 7.030000000e-07 V_low
+ 7.030010000e-07 V_low
+ 7.031000000e-07 V_low
+ 7.031010000e-07 V_low
+ 7.032000000e-07 V_low
+ 7.032010000e-07 V_low
+ 7.033000000e-07 V_low
+ 7.033010000e-07 V_low
+ 7.034000000e-07 V_low
+ 7.034010000e-07 V_low
+ 7.035000000e-07 V_low
+ 7.035010000e-07 V_low
+ 7.036000000e-07 V_low
+ 7.036010000e-07 V_low
+ 7.037000000e-07 V_low
+ 7.037010000e-07 V_low
+ 7.038000000e-07 V_low
+ 7.038010000e-07 V_low
+ 7.039000000e-07 V_low
+ 7.039010000e-07 V_hig
+ 7.040000000e-07 V_hig
+ 7.040010000e-07 V_hig
+ 7.041000000e-07 V_hig
+ 7.041010000e-07 V_hig
+ 7.042000000e-07 V_hig
+ 7.042010000e-07 V_hig
+ 7.043000000e-07 V_hig
+ 7.043010000e-07 V_hig
+ 7.044000000e-07 V_hig
+ 7.044010000e-07 V_hig
+ 7.045000000e-07 V_hig
+ 7.045010000e-07 V_hig
+ 7.046000000e-07 V_hig
+ 7.046010000e-07 V_hig
+ 7.047000000e-07 V_hig
+ 7.047010000e-07 V_hig
+ 7.048000000e-07 V_hig
+ 7.048010000e-07 V_hig
+ 7.049000000e-07 V_hig
+ 7.049010000e-07 V_hig
+ 7.050000000e-07 V_hig
+ 7.050010000e-07 V_hig
+ 7.051000000e-07 V_hig
+ 7.051010000e-07 V_hig
+ 7.052000000e-07 V_hig
+ 7.052010000e-07 V_hig
+ 7.053000000e-07 V_hig
+ 7.053010000e-07 V_hig
+ 7.054000000e-07 V_hig
+ 7.054010000e-07 V_hig
+ 7.055000000e-07 V_hig
+ 7.055010000e-07 V_hig
+ 7.056000000e-07 V_hig
+ 7.056010000e-07 V_hig
+ 7.057000000e-07 V_hig
+ 7.057010000e-07 V_hig
+ 7.058000000e-07 V_hig
+ 7.058010000e-07 V_hig
+ 7.059000000e-07 V_hig
+ 7.059010000e-07 V_low
+ 7.060000000e-07 V_low
+ 7.060010000e-07 V_low
+ 7.061000000e-07 V_low
+ 7.061010000e-07 V_low
+ 7.062000000e-07 V_low
+ 7.062010000e-07 V_low
+ 7.063000000e-07 V_low
+ 7.063010000e-07 V_low
+ 7.064000000e-07 V_low
+ 7.064010000e-07 V_low
+ 7.065000000e-07 V_low
+ 7.065010000e-07 V_low
+ 7.066000000e-07 V_low
+ 7.066010000e-07 V_low
+ 7.067000000e-07 V_low
+ 7.067010000e-07 V_low
+ 7.068000000e-07 V_low
+ 7.068010000e-07 V_low
+ 7.069000000e-07 V_low
+ 7.069010000e-07 V_hig
+ 7.070000000e-07 V_hig
+ 7.070010000e-07 V_hig
+ 7.071000000e-07 V_hig
+ 7.071010000e-07 V_hig
+ 7.072000000e-07 V_hig
+ 7.072010000e-07 V_hig
+ 7.073000000e-07 V_hig
+ 7.073010000e-07 V_hig
+ 7.074000000e-07 V_hig
+ 7.074010000e-07 V_hig
+ 7.075000000e-07 V_hig
+ 7.075010000e-07 V_hig
+ 7.076000000e-07 V_hig
+ 7.076010000e-07 V_hig
+ 7.077000000e-07 V_hig
+ 7.077010000e-07 V_hig
+ 7.078000000e-07 V_hig
+ 7.078010000e-07 V_hig
+ 7.079000000e-07 V_hig
+ 7.079010000e-07 V_low
+ 7.080000000e-07 V_low
+ 7.080010000e-07 V_low
+ 7.081000000e-07 V_low
+ 7.081010000e-07 V_low
+ 7.082000000e-07 V_low
+ 7.082010000e-07 V_low
+ 7.083000000e-07 V_low
+ 7.083010000e-07 V_low
+ 7.084000000e-07 V_low
+ 7.084010000e-07 V_low
+ 7.085000000e-07 V_low
+ 7.085010000e-07 V_low
+ 7.086000000e-07 V_low
+ 7.086010000e-07 V_low
+ 7.087000000e-07 V_low
+ 7.087010000e-07 V_low
+ 7.088000000e-07 V_low
+ 7.088010000e-07 V_low
+ 7.089000000e-07 V_low
+ 7.089010000e-07 V_low
+ 7.090000000e-07 V_low
+ 7.090010000e-07 V_low
+ 7.091000000e-07 V_low
+ 7.091010000e-07 V_low
+ 7.092000000e-07 V_low
+ 7.092010000e-07 V_low
+ 7.093000000e-07 V_low
+ 7.093010000e-07 V_low
+ 7.094000000e-07 V_low
+ 7.094010000e-07 V_low
+ 7.095000000e-07 V_low
+ 7.095010000e-07 V_low
+ 7.096000000e-07 V_low
+ 7.096010000e-07 V_low
+ 7.097000000e-07 V_low
+ 7.097010000e-07 V_low
+ 7.098000000e-07 V_low
+ 7.098010000e-07 V_low
+ 7.099000000e-07 V_low
+ 7.099010000e-07 V_hig
+ 7.100000000e-07 V_hig
+ 7.100010000e-07 V_hig
+ 7.101000000e-07 V_hig
+ 7.101010000e-07 V_hig
+ 7.102000000e-07 V_hig
+ 7.102010000e-07 V_hig
+ 7.103000000e-07 V_hig
+ 7.103010000e-07 V_hig
+ 7.104000000e-07 V_hig
+ 7.104010000e-07 V_hig
+ 7.105000000e-07 V_hig
+ 7.105010000e-07 V_hig
+ 7.106000000e-07 V_hig
+ 7.106010000e-07 V_hig
+ 7.107000000e-07 V_hig
+ 7.107010000e-07 V_hig
+ 7.108000000e-07 V_hig
+ 7.108010000e-07 V_hig
+ 7.109000000e-07 V_hig
+ 7.109010000e-07 V_low
+ 7.110000000e-07 V_low
+ 7.110010000e-07 V_low
+ 7.111000000e-07 V_low
+ 7.111010000e-07 V_low
+ 7.112000000e-07 V_low
+ 7.112010000e-07 V_low
+ 7.113000000e-07 V_low
+ 7.113010000e-07 V_low
+ 7.114000000e-07 V_low
+ 7.114010000e-07 V_low
+ 7.115000000e-07 V_low
+ 7.115010000e-07 V_low
+ 7.116000000e-07 V_low
+ 7.116010000e-07 V_low
+ 7.117000000e-07 V_low
+ 7.117010000e-07 V_low
+ 7.118000000e-07 V_low
+ 7.118010000e-07 V_low
+ 7.119000000e-07 V_low
+ 7.119010000e-07 V_hig
+ 7.120000000e-07 V_hig
+ 7.120010000e-07 V_hig
+ 7.121000000e-07 V_hig
+ 7.121010000e-07 V_hig
+ 7.122000000e-07 V_hig
+ 7.122010000e-07 V_hig
+ 7.123000000e-07 V_hig
+ 7.123010000e-07 V_hig
+ 7.124000000e-07 V_hig
+ 7.124010000e-07 V_hig
+ 7.125000000e-07 V_hig
+ 7.125010000e-07 V_hig
+ 7.126000000e-07 V_hig
+ 7.126010000e-07 V_hig
+ 7.127000000e-07 V_hig
+ 7.127010000e-07 V_hig
+ 7.128000000e-07 V_hig
+ 7.128010000e-07 V_hig
+ 7.129000000e-07 V_hig
+ 7.129010000e-07 V_hig
+ 7.130000000e-07 V_hig
+ 7.130010000e-07 V_hig
+ 7.131000000e-07 V_hig
+ 7.131010000e-07 V_hig
+ 7.132000000e-07 V_hig
+ 7.132010000e-07 V_hig
+ 7.133000000e-07 V_hig
+ 7.133010000e-07 V_hig
+ 7.134000000e-07 V_hig
+ 7.134010000e-07 V_hig
+ 7.135000000e-07 V_hig
+ 7.135010000e-07 V_hig
+ 7.136000000e-07 V_hig
+ 7.136010000e-07 V_hig
+ 7.137000000e-07 V_hig
+ 7.137010000e-07 V_hig
+ 7.138000000e-07 V_hig
+ 7.138010000e-07 V_hig
+ 7.139000000e-07 V_hig
+ 7.139010000e-07 V_hig
+ 7.140000000e-07 V_hig
+ 7.140010000e-07 V_hig
+ 7.141000000e-07 V_hig
+ 7.141010000e-07 V_hig
+ 7.142000000e-07 V_hig
+ 7.142010000e-07 V_hig
+ 7.143000000e-07 V_hig
+ 7.143010000e-07 V_hig
+ 7.144000000e-07 V_hig
+ 7.144010000e-07 V_hig
+ 7.145000000e-07 V_hig
+ 7.145010000e-07 V_hig
+ 7.146000000e-07 V_hig
+ 7.146010000e-07 V_hig
+ 7.147000000e-07 V_hig
+ 7.147010000e-07 V_hig
+ 7.148000000e-07 V_hig
+ 7.148010000e-07 V_hig
+ 7.149000000e-07 V_hig
+ 7.149010000e-07 V_hig
+ 7.150000000e-07 V_hig
+ 7.150010000e-07 V_hig
+ 7.151000000e-07 V_hig
+ 7.151010000e-07 V_hig
+ 7.152000000e-07 V_hig
+ 7.152010000e-07 V_hig
+ 7.153000000e-07 V_hig
+ 7.153010000e-07 V_hig
+ 7.154000000e-07 V_hig
+ 7.154010000e-07 V_hig
+ 7.155000000e-07 V_hig
+ 7.155010000e-07 V_hig
+ 7.156000000e-07 V_hig
+ 7.156010000e-07 V_hig
+ 7.157000000e-07 V_hig
+ 7.157010000e-07 V_hig
+ 7.158000000e-07 V_hig
+ 7.158010000e-07 V_hig
+ 7.159000000e-07 V_hig
+ 7.159010000e-07 V_low
+ 7.160000000e-07 V_low
+ 7.160010000e-07 V_low
+ 7.161000000e-07 V_low
+ 7.161010000e-07 V_low
+ 7.162000000e-07 V_low
+ 7.162010000e-07 V_low
+ 7.163000000e-07 V_low
+ 7.163010000e-07 V_low
+ 7.164000000e-07 V_low
+ 7.164010000e-07 V_low
+ 7.165000000e-07 V_low
+ 7.165010000e-07 V_low
+ 7.166000000e-07 V_low
+ 7.166010000e-07 V_low
+ 7.167000000e-07 V_low
+ 7.167010000e-07 V_low
+ 7.168000000e-07 V_low
+ 7.168010000e-07 V_low
+ 7.169000000e-07 V_low
+ 7.169010000e-07 V_hig
+ 7.170000000e-07 V_hig
+ 7.170010000e-07 V_hig
+ 7.171000000e-07 V_hig
+ 7.171010000e-07 V_hig
+ 7.172000000e-07 V_hig
+ 7.172010000e-07 V_hig
+ 7.173000000e-07 V_hig
+ 7.173010000e-07 V_hig
+ 7.174000000e-07 V_hig
+ 7.174010000e-07 V_hig
+ 7.175000000e-07 V_hig
+ 7.175010000e-07 V_hig
+ 7.176000000e-07 V_hig
+ 7.176010000e-07 V_hig
+ 7.177000000e-07 V_hig
+ 7.177010000e-07 V_hig
+ 7.178000000e-07 V_hig
+ 7.178010000e-07 V_hig
+ 7.179000000e-07 V_hig
+ 7.179010000e-07 V_low
+ 7.180000000e-07 V_low
+ 7.180010000e-07 V_low
+ 7.181000000e-07 V_low
+ 7.181010000e-07 V_low
+ 7.182000000e-07 V_low
+ 7.182010000e-07 V_low
+ 7.183000000e-07 V_low
+ 7.183010000e-07 V_low
+ 7.184000000e-07 V_low
+ 7.184010000e-07 V_low
+ 7.185000000e-07 V_low
+ 7.185010000e-07 V_low
+ 7.186000000e-07 V_low
+ 7.186010000e-07 V_low
+ 7.187000000e-07 V_low
+ 7.187010000e-07 V_low
+ 7.188000000e-07 V_low
+ 7.188010000e-07 V_low
+ 7.189000000e-07 V_low
+ 7.189010000e-07 V_low
+ 7.190000000e-07 V_low
+ 7.190010000e-07 V_low
+ 7.191000000e-07 V_low
+ 7.191010000e-07 V_low
+ 7.192000000e-07 V_low
+ 7.192010000e-07 V_low
+ 7.193000000e-07 V_low
+ 7.193010000e-07 V_low
+ 7.194000000e-07 V_low
+ 7.194010000e-07 V_low
+ 7.195000000e-07 V_low
+ 7.195010000e-07 V_low
+ 7.196000000e-07 V_low
+ 7.196010000e-07 V_low
+ 7.197000000e-07 V_low
+ 7.197010000e-07 V_low
+ 7.198000000e-07 V_low
+ 7.198010000e-07 V_low
+ 7.199000000e-07 V_low
+ 7.199010000e-07 V_hig
+ 7.200000000e-07 V_hig
+ 7.200010000e-07 V_hig
+ 7.201000000e-07 V_hig
+ 7.201010000e-07 V_hig
+ 7.202000000e-07 V_hig
+ 7.202010000e-07 V_hig
+ 7.203000000e-07 V_hig
+ 7.203010000e-07 V_hig
+ 7.204000000e-07 V_hig
+ 7.204010000e-07 V_hig
+ 7.205000000e-07 V_hig
+ 7.205010000e-07 V_hig
+ 7.206000000e-07 V_hig
+ 7.206010000e-07 V_hig
+ 7.207000000e-07 V_hig
+ 7.207010000e-07 V_hig
+ 7.208000000e-07 V_hig
+ 7.208010000e-07 V_hig
+ 7.209000000e-07 V_hig
+ 7.209010000e-07 V_low
+ 7.210000000e-07 V_low
+ 7.210010000e-07 V_low
+ 7.211000000e-07 V_low
+ 7.211010000e-07 V_low
+ 7.212000000e-07 V_low
+ 7.212010000e-07 V_low
+ 7.213000000e-07 V_low
+ 7.213010000e-07 V_low
+ 7.214000000e-07 V_low
+ 7.214010000e-07 V_low
+ 7.215000000e-07 V_low
+ 7.215010000e-07 V_low
+ 7.216000000e-07 V_low
+ 7.216010000e-07 V_low
+ 7.217000000e-07 V_low
+ 7.217010000e-07 V_low
+ 7.218000000e-07 V_low
+ 7.218010000e-07 V_low
+ 7.219000000e-07 V_low
+ 7.219010000e-07 V_hig
+ 7.220000000e-07 V_hig
+ 7.220010000e-07 V_hig
+ 7.221000000e-07 V_hig
+ 7.221010000e-07 V_hig
+ 7.222000000e-07 V_hig
+ 7.222010000e-07 V_hig
+ 7.223000000e-07 V_hig
+ 7.223010000e-07 V_hig
+ 7.224000000e-07 V_hig
+ 7.224010000e-07 V_hig
+ 7.225000000e-07 V_hig
+ 7.225010000e-07 V_hig
+ 7.226000000e-07 V_hig
+ 7.226010000e-07 V_hig
+ 7.227000000e-07 V_hig
+ 7.227010000e-07 V_hig
+ 7.228000000e-07 V_hig
+ 7.228010000e-07 V_hig
+ 7.229000000e-07 V_hig
+ 7.229010000e-07 V_low
+ 7.230000000e-07 V_low
+ 7.230010000e-07 V_low
+ 7.231000000e-07 V_low
+ 7.231010000e-07 V_low
+ 7.232000000e-07 V_low
+ 7.232010000e-07 V_low
+ 7.233000000e-07 V_low
+ 7.233010000e-07 V_low
+ 7.234000000e-07 V_low
+ 7.234010000e-07 V_low
+ 7.235000000e-07 V_low
+ 7.235010000e-07 V_low
+ 7.236000000e-07 V_low
+ 7.236010000e-07 V_low
+ 7.237000000e-07 V_low
+ 7.237010000e-07 V_low
+ 7.238000000e-07 V_low
+ 7.238010000e-07 V_low
+ 7.239000000e-07 V_low
+ 7.239010000e-07 V_hig
+ 7.240000000e-07 V_hig
+ 7.240010000e-07 V_hig
+ 7.241000000e-07 V_hig
+ 7.241010000e-07 V_hig
+ 7.242000000e-07 V_hig
+ 7.242010000e-07 V_hig
+ 7.243000000e-07 V_hig
+ 7.243010000e-07 V_hig
+ 7.244000000e-07 V_hig
+ 7.244010000e-07 V_hig
+ 7.245000000e-07 V_hig
+ 7.245010000e-07 V_hig
+ 7.246000000e-07 V_hig
+ 7.246010000e-07 V_hig
+ 7.247000000e-07 V_hig
+ 7.247010000e-07 V_hig
+ 7.248000000e-07 V_hig
+ 7.248010000e-07 V_hig
+ 7.249000000e-07 V_hig
+ 7.249010000e-07 V_low
+ 7.250000000e-07 V_low
+ 7.250010000e-07 V_low
+ 7.251000000e-07 V_low
+ 7.251010000e-07 V_low
+ 7.252000000e-07 V_low
+ 7.252010000e-07 V_low
+ 7.253000000e-07 V_low
+ 7.253010000e-07 V_low
+ 7.254000000e-07 V_low
+ 7.254010000e-07 V_low
+ 7.255000000e-07 V_low
+ 7.255010000e-07 V_low
+ 7.256000000e-07 V_low
+ 7.256010000e-07 V_low
+ 7.257000000e-07 V_low
+ 7.257010000e-07 V_low
+ 7.258000000e-07 V_low
+ 7.258010000e-07 V_low
+ 7.259000000e-07 V_low
+ 7.259010000e-07 V_low
+ 7.260000000e-07 V_low
+ 7.260010000e-07 V_low
+ 7.261000000e-07 V_low
+ 7.261010000e-07 V_low
+ 7.262000000e-07 V_low
+ 7.262010000e-07 V_low
+ 7.263000000e-07 V_low
+ 7.263010000e-07 V_low
+ 7.264000000e-07 V_low
+ 7.264010000e-07 V_low
+ 7.265000000e-07 V_low
+ 7.265010000e-07 V_low
+ 7.266000000e-07 V_low
+ 7.266010000e-07 V_low
+ 7.267000000e-07 V_low
+ 7.267010000e-07 V_low
+ 7.268000000e-07 V_low
+ 7.268010000e-07 V_low
+ 7.269000000e-07 V_low
+ 7.269010000e-07 V_low
+ 7.270000000e-07 V_low
+ 7.270010000e-07 V_low
+ 7.271000000e-07 V_low
+ 7.271010000e-07 V_low
+ 7.272000000e-07 V_low
+ 7.272010000e-07 V_low
+ 7.273000000e-07 V_low
+ 7.273010000e-07 V_low
+ 7.274000000e-07 V_low
+ 7.274010000e-07 V_low
+ 7.275000000e-07 V_low
+ 7.275010000e-07 V_low
+ 7.276000000e-07 V_low
+ 7.276010000e-07 V_low
+ 7.277000000e-07 V_low
+ 7.277010000e-07 V_low
+ 7.278000000e-07 V_low
+ 7.278010000e-07 V_low
+ 7.279000000e-07 V_low
+ 7.279010000e-07 V_low
+ 7.280000000e-07 V_low
+ 7.280010000e-07 V_low
+ 7.281000000e-07 V_low
+ 7.281010000e-07 V_low
+ 7.282000000e-07 V_low
+ 7.282010000e-07 V_low
+ 7.283000000e-07 V_low
+ 7.283010000e-07 V_low
+ 7.284000000e-07 V_low
+ 7.284010000e-07 V_low
+ 7.285000000e-07 V_low
+ 7.285010000e-07 V_low
+ 7.286000000e-07 V_low
+ 7.286010000e-07 V_low
+ 7.287000000e-07 V_low
+ 7.287010000e-07 V_low
+ 7.288000000e-07 V_low
+ 7.288010000e-07 V_low
+ 7.289000000e-07 V_low
+ 7.289010000e-07 V_low
+ 7.290000000e-07 V_low
+ 7.290010000e-07 V_low
+ 7.291000000e-07 V_low
+ 7.291010000e-07 V_low
+ 7.292000000e-07 V_low
+ 7.292010000e-07 V_low
+ 7.293000000e-07 V_low
+ 7.293010000e-07 V_low
+ 7.294000000e-07 V_low
+ 7.294010000e-07 V_low
+ 7.295000000e-07 V_low
+ 7.295010000e-07 V_low
+ 7.296000000e-07 V_low
+ 7.296010000e-07 V_low
+ 7.297000000e-07 V_low
+ 7.297010000e-07 V_low
+ 7.298000000e-07 V_low
+ 7.298010000e-07 V_low
+ 7.299000000e-07 V_low
+ 7.299010000e-07 V_hig
+ 7.300000000e-07 V_hig
+ 7.300010000e-07 V_hig
+ 7.301000000e-07 V_hig
+ 7.301010000e-07 V_hig
+ 7.302000000e-07 V_hig
+ 7.302010000e-07 V_hig
+ 7.303000000e-07 V_hig
+ 7.303010000e-07 V_hig
+ 7.304000000e-07 V_hig
+ 7.304010000e-07 V_hig
+ 7.305000000e-07 V_hig
+ 7.305010000e-07 V_hig
+ 7.306000000e-07 V_hig
+ 7.306010000e-07 V_hig
+ 7.307000000e-07 V_hig
+ 7.307010000e-07 V_hig
+ 7.308000000e-07 V_hig
+ 7.308010000e-07 V_hig
+ 7.309000000e-07 V_hig
+ 7.309010000e-07 V_low
+ 7.310000000e-07 V_low
+ 7.310010000e-07 V_low
+ 7.311000000e-07 V_low
+ 7.311010000e-07 V_low
+ 7.312000000e-07 V_low
+ 7.312010000e-07 V_low
+ 7.313000000e-07 V_low
+ 7.313010000e-07 V_low
+ 7.314000000e-07 V_low
+ 7.314010000e-07 V_low
+ 7.315000000e-07 V_low
+ 7.315010000e-07 V_low
+ 7.316000000e-07 V_low
+ 7.316010000e-07 V_low
+ 7.317000000e-07 V_low
+ 7.317010000e-07 V_low
+ 7.318000000e-07 V_low
+ 7.318010000e-07 V_low
+ 7.319000000e-07 V_low
+ 7.319010000e-07 V_hig
+ 7.320000000e-07 V_hig
+ 7.320010000e-07 V_hig
+ 7.321000000e-07 V_hig
+ 7.321010000e-07 V_hig
+ 7.322000000e-07 V_hig
+ 7.322010000e-07 V_hig
+ 7.323000000e-07 V_hig
+ 7.323010000e-07 V_hig
+ 7.324000000e-07 V_hig
+ 7.324010000e-07 V_hig
+ 7.325000000e-07 V_hig
+ 7.325010000e-07 V_hig
+ 7.326000000e-07 V_hig
+ 7.326010000e-07 V_hig
+ 7.327000000e-07 V_hig
+ 7.327010000e-07 V_hig
+ 7.328000000e-07 V_hig
+ 7.328010000e-07 V_hig
+ 7.329000000e-07 V_hig
+ 7.329010000e-07 V_hig
+ 7.330000000e-07 V_hig
+ 7.330010000e-07 V_hig
+ 7.331000000e-07 V_hig
+ 7.331010000e-07 V_hig
+ 7.332000000e-07 V_hig
+ 7.332010000e-07 V_hig
+ 7.333000000e-07 V_hig
+ 7.333010000e-07 V_hig
+ 7.334000000e-07 V_hig
+ 7.334010000e-07 V_hig
+ 7.335000000e-07 V_hig
+ 7.335010000e-07 V_hig
+ 7.336000000e-07 V_hig
+ 7.336010000e-07 V_hig
+ 7.337000000e-07 V_hig
+ 7.337010000e-07 V_hig
+ 7.338000000e-07 V_hig
+ 7.338010000e-07 V_hig
+ 7.339000000e-07 V_hig
+ 7.339010000e-07 V_low
+ 7.340000000e-07 V_low
+ 7.340010000e-07 V_low
+ 7.341000000e-07 V_low
+ 7.341010000e-07 V_low
+ 7.342000000e-07 V_low
+ 7.342010000e-07 V_low
+ 7.343000000e-07 V_low
+ 7.343010000e-07 V_low
+ 7.344000000e-07 V_low
+ 7.344010000e-07 V_low
+ 7.345000000e-07 V_low
+ 7.345010000e-07 V_low
+ 7.346000000e-07 V_low
+ 7.346010000e-07 V_low
+ 7.347000000e-07 V_low
+ 7.347010000e-07 V_low
+ 7.348000000e-07 V_low
+ 7.348010000e-07 V_low
+ 7.349000000e-07 V_low
+ 7.349010000e-07 V_low
+ 7.350000000e-07 V_low
+ 7.350010000e-07 V_low
+ 7.351000000e-07 V_low
+ 7.351010000e-07 V_low
+ 7.352000000e-07 V_low
+ 7.352010000e-07 V_low
+ 7.353000000e-07 V_low
+ 7.353010000e-07 V_low
+ 7.354000000e-07 V_low
+ 7.354010000e-07 V_low
+ 7.355000000e-07 V_low
+ 7.355010000e-07 V_low
+ 7.356000000e-07 V_low
+ 7.356010000e-07 V_low
+ 7.357000000e-07 V_low
+ 7.357010000e-07 V_low
+ 7.358000000e-07 V_low
+ 7.358010000e-07 V_low
+ 7.359000000e-07 V_low
+ 7.359010000e-07 V_hig
+ 7.360000000e-07 V_hig
+ 7.360010000e-07 V_hig
+ 7.361000000e-07 V_hig
+ 7.361010000e-07 V_hig
+ 7.362000000e-07 V_hig
+ 7.362010000e-07 V_hig
+ 7.363000000e-07 V_hig
+ 7.363010000e-07 V_hig
+ 7.364000000e-07 V_hig
+ 7.364010000e-07 V_hig
+ 7.365000000e-07 V_hig
+ 7.365010000e-07 V_hig
+ 7.366000000e-07 V_hig
+ 7.366010000e-07 V_hig
+ 7.367000000e-07 V_hig
+ 7.367010000e-07 V_hig
+ 7.368000000e-07 V_hig
+ 7.368010000e-07 V_hig
+ 7.369000000e-07 V_hig
+ 7.369010000e-07 V_low
+ 7.370000000e-07 V_low
+ 7.370010000e-07 V_low
+ 7.371000000e-07 V_low
+ 7.371010000e-07 V_low
+ 7.372000000e-07 V_low
+ 7.372010000e-07 V_low
+ 7.373000000e-07 V_low
+ 7.373010000e-07 V_low
+ 7.374000000e-07 V_low
+ 7.374010000e-07 V_low
+ 7.375000000e-07 V_low
+ 7.375010000e-07 V_low
+ 7.376000000e-07 V_low
+ 7.376010000e-07 V_low
+ 7.377000000e-07 V_low
+ 7.377010000e-07 V_low
+ 7.378000000e-07 V_low
+ 7.378010000e-07 V_low
+ 7.379000000e-07 V_low
+ 7.379010000e-07 V_hig
+ 7.380000000e-07 V_hig
+ 7.380010000e-07 V_hig
+ 7.381000000e-07 V_hig
+ 7.381010000e-07 V_hig
+ 7.382000000e-07 V_hig
+ 7.382010000e-07 V_hig
+ 7.383000000e-07 V_hig
+ 7.383010000e-07 V_hig
+ 7.384000000e-07 V_hig
+ 7.384010000e-07 V_hig
+ 7.385000000e-07 V_hig
+ 7.385010000e-07 V_hig
+ 7.386000000e-07 V_hig
+ 7.386010000e-07 V_hig
+ 7.387000000e-07 V_hig
+ 7.387010000e-07 V_hig
+ 7.388000000e-07 V_hig
+ 7.388010000e-07 V_hig
+ 7.389000000e-07 V_hig
+ 7.389010000e-07 V_low
+ 7.390000000e-07 V_low
+ 7.390010000e-07 V_low
+ 7.391000000e-07 V_low
+ 7.391010000e-07 V_low
+ 7.392000000e-07 V_low
+ 7.392010000e-07 V_low
+ 7.393000000e-07 V_low
+ 7.393010000e-07 V_low
+ 7.394000000e-07 V_low
+ 7.394010000e-07 V_low
+ 7.395000000e-07 V_low
+ 7.395010000e-07 V_low
+ 7.396000000e-07 V_low
+ 7.396010000e-07 V_low
+ 7.397000000e-07 V_low
+ 7.397010000e-07 V_low
+ 7.398000000e-07 V_low
+ 7.398010000e-07 V_low
+ 7.399000000e-07 V_low
+ 7.399010000e-07 V_hig
+ 7.400000000e-07 V_hig
+ 7.400010000e-07 V_hig
+ 7.401000000e-07 V_hig
+ 7.401010000e-07 V_hig
+ 7.402000000e-07 V_hig
+ 7.402010000e-07 V_hig
+ 7.403000000e-07 V_hig
+ 7.403010000e-07 V_hig
+ 7.404000000e-07 V_hig
+ 7.404010000e-07 V_hig
+ 7.405000000e-07 V_hig
+ 7.405010000e-07 V_hig
+ 7.406000000e-07 V_hig
+ 7.406010000e-07 V_hig
+ 7.407000000e-07 V_hig
+ 7.407010000e-07 V_hig
+ 7.408000000e-07 V_hig
+ 7.408010000e-07 V_hig
+ 7.409000000e-07 V_hig
+ 7.409010000e-07 V_low
+ 7.410000000e-07 V_low
+ 7.410010000e-07 V_low
+ 7.411000000e-07 V_low
+ 7.411010000e-07 V_low
+ 7.412000000e-07 V_low
+ 7.412010000e-07 V_low
+ 7.413000000e-07 V_low
+ 7.413010000e-07 V_low
+ 7.414000000e-07 V_low
+ 7.414010000e-07 V_low
+ 7.415000000e-07 V_low
+ 7.415010000e-07 V_low
+ 7.416000000e-07 V_low
+ 7.416010000e-07 V_low
+ 7.417000000e-07 V_low
+ 7.417010000e-07 V_low
+ 7.418000000e-07 V_low
+ 7.418010000e-07 V_low
+ 7.419000000e-07 V_low
+ 7.419010000e-07 V_hig
+ 7.420000000e-07 V_hig
+ 7.420010000e-07 V_hig
+ 7.421000000e-07 V_hig
+ 7.421010000e-07 V_hig
+ 7.422000000e-07 V_hig
+ 7.422010000e-07 V_hig
+ 7.423000000e-07 V_hig
+ 7.423010000e-07 V_hig
+ 7.424000000e-07 V_hig
+ 7.424010000e-07 V_hig
+ 7.425000000e-07 V_hig
+ 7.425010000e-07 V_hig
+ 7.426000000e-07 V_hig
+ 7.426010000e-07 V_hig
+ 7.427000000e-07 V_hig
+ 7.427010000e-07 V_hig
+ 7.428000000e-07 V_hig
+ 7.428010000e-07 V_hig
+ 7.429000000e-07 V_hig
+ 7.429010000e-07 V_low
+ 7.430000000e-07 V_low
+ 7.430010000e-07 V_low
+ 7.431000000e-07 V_low
+ 7.431010000e-07 V_low
+ 7.432000000e-07 V_low
+ 7.432010000e-07 V_low
+ 7.433000000e-07 V_low
+ 7.433010000e-07 V_low
+ 7.434000000e-07 V_low
+ 7.434010000e-07 V_low
+ 7.435000000e-07 V_low
+ 7.435010000e-07 V_low
+ 7.436000000e-07 V_low
+ 7.436010000e-07 V_low
+ 7.437000000e-07 V_low
+ 7.437010000e-07 V_low
+ 7.438000000e-07 V_low
+ 7.438010000e-07 V_low
+ 7.439000000e-07 V_low
+ 7.439010000e-07 V_low
+ 7.440000000e-07 V_low
+ 7.440010000e-07 V_low
+ 7.441000000e-07 V_low
+ 7.441010000e-07 V_low
+ 7.442000000e-07 V_low
+ 7.442010000e-07 V_low
+ 7.443000000e-07 V_low
+ 7.443010000e-07 V_low
+ 7.444000000e-07 V_low
+ 7.444010000e-07 V_low
+ 7.445000000e-07 V_low
+ 7.445010000e-07 V_low
+ 7.446000000e-07 V_low
+ 7.446010000e-07 V_low
+ 7.447000000e-07 V_low
+ 7.447010000e-07 V_low
+ 7.448000000e-07 V_low
+ 7.448010000e-07 V_low
+ 7.449000000e-07 V_low
+ 7.449010000e-07 V_low
+ 7.450000000e-07 V_low
+ 7.450010000e-07 V_low
+ 7.451000000e-07 V_low
+ 7.451010000e-07 V_low
+ 7.452000000e-07 V_low
+ 7.452010000e-07 V_low
+ 7.453000000e-07 V_low
+ 7.453010000e-07 V_low
+ 7.454000000e-07 V_low
+ 7.454010000e-07 V_low
+ 7.455000000e-07 V_low
+ 7.455010000e-07 V_low
+ 7.456000000e-07 V_low
+ 7.456010000e-07 V_low
+ 7.457000000e-07 V_low
+ 7.457010000e-07 V_low
+ 7.458000000e-07 V_low
+ 7.458010000e-07 V_low
+ 7.459000000e-07 V_low
+ 7.459010000e-07 V_low
+ 7.460000000e-07 V_low
+ 7.460010000e-07 V_low
+ 7.461000000e-07 V_low
+ 7.461010000e-07 V_low
+ 7.462000000e-07 V_low
+ 7.462010000e-07 V_low
+ 7.463000000e-07 V_low
+ 7.463010000e-07 V_low
+ 7.464000000e-07 V_low
+ 7.464010000e-07 V_low
+ 7.465000000e-07 V_low
+ 7.465010000e-07 V_low
+ 7.466000000e-07 V_low
+ 7.466010000e-07 V_low
+ 7.467000000e-07 V_low
+ 7.467010000e-07 V_low
+ 7.468000000e-07 V_low
+ 7.468010000e-07 V_low
+ 7.469000000e-07 V_low
+ 7.469010000e-07 V_hig
+ 7.470000000e-07 V_hig
+ 7.470010000e-07 V_hig
+ 7.471000000e-07 V_hig
+ 7.471010000e-07 V_hig
+ 7.472000000e-07 V_hig
+ 7.472010000e-07 V_hig
+ 7.473000000e-07 V_hig
+ 7.473010000e-07 V_hig
+ 7.474000000e-07 V_hig
+ 7.474010000e-07 V_hig
+ 7.475000000e-07 V_hig
+ 7.475010000e-07 V_hig
+ 7.476000000e-07 V_hig
+ 7.476010000e-07 V_hig
+ 7.477000000e-07 V_hig
+ 7.477010000e-07 V_hig
+ 7.478000000e-07 V_hig
+ 7.478010000e-07 V_hig
+ 7.479000000e-07 V_hig
+ 7.479010000e-07 V_low
+ 7.480000000e-07 V_low
+ 7.480010000e-07 V_low
+ 7.481000000e-07 V_low
+ 7.481010000e-07 V_low
+ 7.482000000e-07 V_low
+ 7.482010000e-07 V_low
+ 7.483000000e-07 V_low
+ 7.483010000e-07 V_low
+ 7.484000000e-07 V_low
+ 7.484010000e-07 V_low
+ 7.485000000e-07 V_low
+ 7.485010000e-07 V_low
+ 7.486000000e-07 V_low
+ 7.486010000e-07 V_low
+ 7.487000000e-07 V_low
+ 7.487010000e-07 V_low
+ 7.488000000e-07 V_low
+ 7.488010000e-07 V_low
+ 7.489000000e-07 V_low
+ 7.489010000e-07 V_low
+ 7.490000000e-07 V_low
+ 7.490010000e-07 V_low
+ 7.491000000e-07 V_low
+ 7.491010000e-07 V_low
+ 7.492000000e-07 V_low
+ 7.492010000e-07 V_low
+ 7.493000000e-07 V_low
+ 7.493010000e-07 V_low
+ 7.494000000e-07 V_low
+ 7.494010000e-07 V_low
+ 7.495000000e-07 V_low
+ 7.495010000e-07 V_low
+ 7.496000000e-07 V_low
+ 7.496010000e-07 V_low
+ 7.497000000e-07 V_low
+ 7.497010000e-07 V_low
+ 7.498000000e-07 V_low
+ 7.498010000e-07 V_low
+ 7.499000000e-07 V_low
+ 7.499010000e-07 V_hig
+ 7.500000000e-07 V_hig
+ 7.500010000e-07 V_hig
+ 7.501000000e-07 V_hig
+ 7.501010000e-07 V_hig
+ 7.502000000e-07 V_hig
+ 7.502010000e-07 V_hig
+ 7.503000000e-07 V_hig
+ 7.503010000e-07 V_hig
+ 7.504000000e-07 V_hig
+ 7.504010000e-07 V_hig
+ 7.505000000e-07 V_hig
+ 7.505010000e-07 V_hig
+ 7.506000000e-07 V_hig
+ 7.506010000e-07 V_hig
+ 7.507000000e-07 V_hig
+ 7.507010000e-07 V_hig
+ 7.508000000e-07 V_hig
+ 7.508010000e-07 V_hig
+ 7.509000000e-07 V_hig
+ 7.509010000e-07 V_low
+ 7.510000000e-07 V_low
+ 7.510010000e-07 V_low
+ 7.511000000e-07 V_low
+ 7.511010000e-07 V_low
+ 7.512000000e-07 V_low
+ 7.512010000e-07 V_low
+ 7.513000000e-07 V_low
+ 7.513010000e-07 V_low
+ 7.514000000e-07 V_low
+ 7.514010000e-07 V_low
+ 7.515000000e-07 V_low
+ 7.515010000e-07 V_low
+ 7.516000000e-07 V_low
+ 7.516010000e-07 V_low
+ 7.517000000e-07 V_low
+ 7.517010000e-07 V_low
+ 7.518000000e-07 V_low
+ 7.518010000e-07 V_low
+ 7.519000000e-07 V_low
+ 7.519010000e-07 V_hig
+ 7.520000000e-07 V_hig
+ 7.520010000e-07 V_hig
+ 7.521000000e-07 V_hig
+ 7.521010000e-07 V_hig
+ 7.522000000e-07 V_hig
+ 7.522010000e-07 V_hig
+ 7.523000000e-07 V_hig
+ 7.523010000e-07 V_hig
+ 7.524000000e-07 V_hig
+ 7.524010000e-07 V_hig
+ 7.525000000e-07 V_hig
+ 7.525010000e-07 V_hig
+ 7.526000000e-07 V_hig
+ 7.526010000e-07 V_hig
+ 7.527000000e-07 V_hig
+ 7.527010000e-07 V_hig
+ 7.528000000e-07 V_hig
+ 7.528010000e-07 V_hig
+ 7.529000000e-07 V_hig
+ 7.529010000e-07 V_hig
+ 7.530000000e-07 V_hig
+ 7.530010000e-07 V_hig
+ 7.531000000e-07 V_hig
+ 7.531010000e-07 V_hig
+ 7.532000000e-07 V_hig
+ 7.532010000e-07 V_hig
+ 7.533000000e-07 V_hig
+ 7.533010000e-07 V_hig
+ 7.534000000e-07 V_hig
+ 7.534010000e-07 V_hig
+ 7.535000000e-07 V_hig
+ 7.535010000e-07 V_hig
+ 7.536000000e-07 V_hig
+ 7.536010000e-07 V_hig
+ 7.537000000e-07 V_hig
+ 7.537010000e-07 V_hig
+ 7.538000000e-07 V_hig
+ 7.538010000e-07 V_hig
+ 7.539000000e-07 V_hig
+ 7.539010000e-07 V_low
+ 7.540000000e-07 V_low
+ 7.540010000e-07 V_low
+ 7.541000000e-07 V_low
+ 7.541010000e-07 V_low
+ 7.542000000e-07 V_low
+ 7.542010000e-07 V_low
+ 7.543000000e-07 V_low
+ 7.543010000e-07 V_low
+ 7.544000000e-07 V_low
+ 7.544010000e-07 V_low
+ 7.545000000e-07 V_low
+ 7.545010000e-07 V_low
+ 7.546000000e-07 V_low
+ 7.546010000e-07 V_low
+ 7.547000000e-07 V_low
+ 7.547010000e-07 V_low
+ 7.548000000e-07 V_low
+ 7.548010000e-07 V_low
+ 7.549000000e-07 V_low
+ 7.549010000e-07 V_low
+ 7.550000000e-07 V_low
+ 7.550010000e-07 V_low
+ 7.551000000e-07 V_low
+ 7.551010000e-07 V_low
+ 7.552000000e-07 V_low
+ 7.552010000e-07 V_low
+ 7.553000000e-07 V_low
+ 7.553010000e-07 V_low
+ 7.554000000e-07 V_low
+ 7.554010000e-07 V_low
+ 7.555000000e-07 V_low
+ 7.555010000e-07 V_low
+ 7.556000000e-07 V_low
+ 7.556010000e-07 V_low
+ 7.557000000e-07 V_low
+ 7.557010000e-07 V_low
+ 7.558000000e-07 V_low
+ 7.558010000e-07 V_low
+ 7.559000000e-07 V_low
+ 7.559010000e-07 V_hig
+ 7.560000000e-07 V_hig
+ 7.560010000e-07 V_hig
+ 7.561000000e-07 V_hig
+ 7.561010000e-07 V_hig
+ 7.562000000e-07 V_hig
+ 7.562010000e-07 V_hig
+ 7.563000000e-07 V_hig
+ 7.563010000e-07 V_hig
+ 7.564000000e-07 V_hig
+ 7.564010000e-07 V_hig
+ 7.565000000e-07 V_hig
+ 7.565010000e-07 V_hig
+ 7.566000000e-07 V_hig
+ 7.566010000e-07 V_hig
+ 7.567000000e-07 V_hig
+ 7.567010000e-07 V_hig
+ 7.568000000e-07 V_hig
+ 7.568010000e-07 V_hig
+ 7.569000000e-07 V_hig
+ 7.569010000e-07 V_hig
+ 7.570000000e-07 V_hig
+ 7.570010000e-07 V_hig
+ 7.571000000e-07 V_hig
+ 7.571010000e-07 V_hig
+ 7.572000000e-07 V_hig
+ 7.572010000e-07 V_hig
+ 7.573000000e-07 V_hig
+ 7.573010000e-07 V_hig
+ 7.574000000e-07 V_hig
+ 7.574010000e-07 V_hig
+ 7.575000000e-07 V_hig
+ 7.575010000e-07 V_hig
+ 7.576000000e-07 V_hig
+ 7.576010000e-07 V_hig
+ 7.577000000e-07 V_hig
+ 7.577010000e-07 V_hig
+ 7.578000000e-07 V_hig
+ 7.578010000e-07 V_hig
+ 7.579000000e-07 V_hig
+ 7.579010000e-07 V_hig
+ 7.580000000e-07 V_hig
+ 7.580010000e-07 V_hig
+ 7.581000000e-07 V_hig
+ 7.581010000e-07 V_hig
+ 7.582000000e-07 V_hig
+ 7.582010000e-07 V_hig
+ 7.583000000e-07 V_hig
+ 7.583010000e-07 V_hig
+ 7.584000000e-07 V_hig
+ 7.584010000e-07 V_hig
+ 7.585000000e-07 V_hig
+ 7.585010000e-07 V_hig
+ 7.586000000e-07 V_hig
+ 7.586010000e-07 V_hig
+ 7.587000000e-07 V_hig
+ 7.587010000e-07 V_hig
+ 7.588000000e-07 V_hig
+ 7.588010000e-07 V_hig
+ 7.589000000e-07 V_hig
+ 7.589010000e-07 V_low
+ 7.590000000e-07 V_low
+ 7.590010000e-07 V_low
+ 7.591000000e-07 V_low
+ 7.591010000e-07 V_low
+ 7.592000000e-07 V_low
+ 7.592010000e-07 V_low
+ 7.593000000e-07 V_low
+ 7.593010000e-07 V_low
+ 7.594000000e-07 V_low
+ 7.594010000e-07 V_low
+ 7.595000000e-07 V_low
+ 7.595010000e-07 V_low
+ 7.596000000e-07 V_low
+ 7.596010000e-07 V_low
+ 7.597000000e-07 V_low
+ 7.597010000e-07 V_low
+ 7.598000000e-07 V_low
+ 7.598010000e-07 V_low
+ 7.599000000e-07 V_low
+ 7.599010000e-07 V_hig
+ 7.600000000e-07 V_hig
+ 7.600010000e-07 V_hig
+ 7.601000000e-07 V_hig
+ 7.601010000e-07 V_hig
+ 7.602000000e-07 V_hig
+ 7.602010000e-07 V_hig
+ 7.603000000e-07 V_hig
+ 7.603010000e-07 V_hig
+ 7.604000000e-07 V_hig
+ 7.604010000e-07 V_hig
+ 7.605000000e-07 V_hig
+ 7.605010000e-07 V_hig
+ 7.606000000e-07 V_hig
+ 7.606010000e-07 V_hig
+ 7.607000000e-07 V_hig
+ 7.607010000e-07 V_hig
+ 7.608000000e-07 V_hig
+ 7.608010000e-07 V_hig
+ 7.609000000e-07 V_hig
+ 7.609010000e-07 V_low
+ 7.610000000e-07 V_low
+ 7.610010000e-07 V_low
+ 7.611000000e-07 V_low
+ 7.611010000e-07 V_low
+ 7.612000000e-07 V_low
+ 7.612010000e-07 V_low
+ 7.613000000e-07 V_low
+ 7.613010000e-07 V_low
+ 7.614000000e-07 V_low
+ 7.614010000e-07 V_low
+ 7.615000000e-07 V_low
+ 7.615010000e-07 V_low
+ 7.616000000e-07 V_low
+ 7.616010000e-07 V_low
+ 7.617000000e-07 V_low
+ 7.617010000e-07 V_low
+ 7.618000000e-07 V_low
+ 7.618010000e-07 V_low
+ 7.619000000e-07 V_low
+ 7.619010000e-07 V_low
+ 7.620000000e-07 V_low
+ 7.620010000e-07 V_low
+ 7.621000000e-07 V_low
+ 7.621010000e-07 V_low
+ 7.622000000e-07 V_low
+ 7.622010000e-07 V_low
+ 7.623000000e-07 V_low
+ 7.623010000e-07 V_low
+ 7.624000000e-07 V_low
+ 7.624010000e-07 V_low
+ 7.625000000e-07 V_low
+ 7.625010000e-07 V_low
+ 7.626000000e-07 V_low
+ 7.626010000e-07 V_low
+ 7.627000000e-07 V_low
+ 7.627010000e-07 V_low
+ 7.628000000e-07 V_low
+ 7.628010000e-07 V_low
+ 7.629000000e-07 V_low
+ 7.629010000e-07 V_low
+ 7.630000000e-07 V_low
+ 7.630010000e-07 V_low
+ 7.631000000e-07 V_low
+ 7.631010000e-07 V_low
+ 7.632000000e-07 V_low
+ 7.632010000e-07 V_low
+ 7.633000000e-07 V_low
+ 7.633010000e-07 V_low
+ 7.634000000e-07 V_low
+ 7.634010000e-07 V_low
+ 7.635000000e-07 V_low
+ 7.635010000e-07 V_low
+ 7.636000000e-07 V_low
+ 7.636010000e-07 V_low
+ 7.637000000e-07 V_low
+ 7.637010000e-07 V_low
+ 7.638000000e-07 V_low
+ 7.638010000e-07 V_low
+ 7.639000000e-07 V_low
+ 7.639010000e-07 V_hig
+ 7.640000000e-07 V_hig
+ 7.640010000e-07 V_hig
+ 7.641000000e-07 V_hig
+ 7.641010000e-07 V_hig
+ 7.642000000e-07 V_hig
+ 7.642010000e-07 V_hig
+ 7.643000000e-07 V_hig
+ 7.643010000e-07 V_hig
+ 7.644000000e-07 V_hig
+ 7.644010000e-07 V_hig
+ 7.645000000e-07 V_hig
+ 7.645010000e-07 V_hig
+ 7.646000000e-07 V_hig
+ 7.646010000e-07 V_hig
+ 7.647000000e-07 V_hig
+ 7.647010000e-07 V_hig
+ 7.648000000e-07 V_hig
+ 7.648010000e-07 V_hig
+ 7.649000000e-07 V_hig
+ 7.649010000e-07 V_hig
+ 7.650000000e-07 V_hig
+ 7.650010000e-07 V_hig
+ 7.651000000e-07 V_hig
+ 7.651010000e-07 V_hig
+ 7.652000000e-07 V_hig
+ 7.652010000e-07 V_hig
+ 7.653000000e-07 V_hig
+ 7.653010000e-07 V_hig
+ 7.654000000e-07 V_hig
+ 7.654010000e-07 V_hig
+ 7.655000000e-07 V_hig
+ 7.655010000e-07 V_hig
+ 7.656000000e-07 V_hig
+ 7.656010000e-07 V_hig
+ 7.657000000e-07 V_hig
+ 7.657010000e-07 V_hig
+ 7.658000000e-07 V_hig
+ 7.658010000e-07 V_hig
+ 7.659000000e-07 V_hig
+ 7.659010000e-07 V_hig
+ 7.660000000e-07 V_hig
+ 7.660010000e-07 V_hig
+ 7.661000000e-07 V_hig
+ 7.661010000e-07 V_hig
+ 7.662000000e-07 V_hig
+ 7.662010000e-07 V_hig
+ 7.663000000e-07 V_hig
+ 7.663010000e-07 V_hig
+ 7.664000000e-07 V_hig
+ 7.664010000e-07 V_hig
+ 7.665000000e-07 V_hig
+ 7.665010000e-07 V_hig
+ 7.666000000e-07 V_hig
+ 7.666010000e-07 V_hig
+ 7.667000000e-07 V_hig
+ 7.667010000e-07 V_hig
+ 7.668000000e-07 V_hig
+ 7.668010000e-07 V_hig
+ 7.669000000e-07 V_hig
+ 7.669010000e-07 V_hig
+ 7.670000000e-07 V_hig
+ 7.670010000e-07 V_hig
+ 7.671000000e-07 V_hig
+ 7.671010000e-07 V_hig
+ 7.672000000e-07 V_hig
+ 7.672010000e-07 V_hig
+ 7.673000000e-07 V_hig
+ 7.673010000e-07 V_hig
+ 7.674000000e-07 V_hig
+ 7.674010000e-07 V_hig
+ 7.675000000e-07 V_hig
+ 7.675010000e-07 V_hig
+ 7.676000000e-07 V_hig
+ 7.676010000e-07 V_hig
+ 7.677000000e-07 V_hig
+ 7.677010000e-07 V_hig
+ 7.678000000e-07 V_hig
+ 7.678010000e-07 V_hig
+ 7.679000000e-07 V_hig
+ 7.679010000e-07 V_low
+ 7.680000000e-07 V_low
+ 7.680010000e-07 V_low
+ 7.681000000e-07 V_low
+ 7.681010000e-07 V_low
+ 7.682000000e-07 V_low
+ 7.682010000e-07 V_low
+ 7.683000000e-07 V_low
+ 7.683010000e-07 V_low
+ 7.684000000e-07 V_low
+ 7.684010000e-07 V_low
+ 7.685000000e-07 V_low
+ 7.685010000e-07 V_low
+ 7.686000000e-07 V_low
+ 7.686010000e-07 V_low
+ 7.687000000e-07 V_low
+ 7.687010000e-07 V_low
+ 7.688000000e-07 V_low
+ 7.688010000e-07 V_low
+ 7.689000000e-07 V_low
+ 7.689010000e-07 V_low
+ 7.690000000e-07 V_low
+ 7.690010000e-07 V_low
+ 7.691000000e-07 V_low
+ 7.691010000e-07 V_low
+ 7.692000000e-07 V_low
+ 7.692010000e-07 V_low
+ 7.693000000e-07 V_low
+ 7.693010000e-07 V_low
+ 7.694000000e-07 V_low
+ 7.694010000e-07 V_low
+ 7.695000000e-07 V_low
+ 7.695010000e-07 V_low
+ 7.696000000e-07 V_low
+ 7.696010000e-07 V_low
+ 7.697000000e-07 V_low
+ 7.697010000e-07 V_low
+ 7.698000000e-07 V_low
+ 7.698010000e-07 V_low
+ 7.699000000e-07 V_low
+ 7.699010000e-07 V_hig
+ 7.700000000e-07 V_hig
+ 7.700010000e-07 V_hig
+ 7.701000000e-07 V_hig
+ 7.701010000e-07 V_hig
+ 7.702000000e-07 V_hig
+ 7.702010000e-07 V_hig
+ 7.703000000e-07 V_hig
+ 7.703010000e-07 V_hig
+ 7.704000000e-07 V_hig
+ 7.704010000e-07 V_hig
+ 7.705000000e-07 V_hig
+ 7.705010000e-07 V_hig
+ 7.706000000e-07 V_hig
+ 7.706010000e-07 V_hig
+ 7.707000000e-07 V_hig
+ 7.707010000e-07 V_hig
+ 7.708000000e-07 V_hig
+ 7.708010000e-07 V_hig
+ 7.709000000e-07 V_hig
+ 7.709010000e-07 V_low
+ 7.710000000e-07 V_low
+ 7.710010000e-07 V_low
+ 7.711000000e-07 V_low
+ 7.711010000e-07 V_low
+ 7.712000000e-07 V_low
+ 7.712010000e-07 V_low
+ 7.713000000e-07 V_low
+ 7.713010000e-07 V_low
+ 7.714000000e-07 V_low
+ 7.714010000e-07 V_low
+ 7.715000000e-07 V_low
+ 7.715010000e-07 V_low
+ 7.716000000e-07 V_low
+ 7.716010000e-07 V_low
+ 7.717000000e-07 V_low
+ 7.717010000e-07 V_low
+ 7.718000000e-07 V_low
+ 7.718010000e-07 V_low
+ 7.719000000e-07 V_low
+ 7.719010000e-07 V_low
+ 7.720000000e-07 V_low
+ 7.720010000e-07 V_low
+ 7.721000000e-07 V_low
+ 7.721010000e-07 V_low
+ 7.722000000e-07 V_low
+ 7.722010000e-07 V_low
+ 7.723000000e-07 V_low
+ 7.723010000e-07 V_low
+ 7.724000000e-07 V_low
+ 7.724010000e-07 V_low
+ 7.725000000e-07 V_low
+ 7.725010000e-07 V_low
+ 7.726000000e-07 V_low
+ 7.726010000e-07 V_low
+ 7.727000000e-07 V_low
+ 7.727010000e-07 V_low
+ 7.728000000e-07 V_low
+ 7.728010000e-07 V_low
+ 7.729000000e-07 V_low
+ 7.729010000e-07 V_hig
+ 7.730000000e-07 V_hig
+ 7.730010000e-07 V_hig
+ 7.731000000e-07 V_hig
+ 7.731010000e-07 V_hig
+ 7.732000000e-07 V_hig
+ 7.732010000e-07 V_hig
+ 7.733000000e-07 V_hig
+ 7.733010000e-07 V_hig
+ 7.734000000e-07 V_hig
+ 7.734010000e-07 V_hig
+ 7.735000000e-07 V_hig
+ 7.735010000e-07 V_hig
+ 7.736000000e-07 V_hig
+ 7.736010000e-07 V_hig
+ 7.737000000e-07 V_hig
+ 7.737010000e-07 V_hig
+ 7.738000000e-07 V_hig
+ 7.738010000e-07 V_hig
+ 7.739000000e-07 V_hig
+ 7.739010000e-07 V_low
+ 7.740000000e-07 V_low
+ 7.740010000e-07 V_low
+ 7.741000000e-07 V_low
+ 7.741010000e-07 V_low
+ 7.742000000e-07 V_low
+ 7.742010000e-07 V_low
+ 7.743000000e-07 V_low
+ 7.743010000e-07 V_low
+ 7.744000000e-07 V_low
+ 7.744010000e-07 V_low
+ 7.745000000e-07 V_low
+ 7.745010000e-07 V_low
+ 7.746000000e-07 V_low
+ 7.746010000e-07 V_low
+ 7.747000000e-07 V_low
+ 7.747010000e-07 V_low
+ 7.748000000e-07 V_low
+ 7.748010000e-07 V_low
+ 7.749000000e-07 V_low
+ 7.749010000e-07 V_low
+ 7.750000000e-07 V_low
+ 7.750010000e-07 V_low
+ 7.751000000e-07 V_low
+ 7.751010000e-07 V_low
+ 7.752000000e-07 V_low
+ 7.752010000e-07 V_low
+ 7.753000000e-07 V_low
+ 7.753010000e-07 V_low
+ 7.754000000e-07 V_low
+ 7.754010000e-07 V_low
+ 7.755000000e-07 V_low
+ 7.755010000e-07 V_low
+ 7.756000000e-07 V_low
+ 7.756010000e-07 V_low
+ 7.757000000e-07 V_low
+ 7.757010000e-07 V_low
+ 7.758000000e-07 V_low
+ 7.758010000e-07 V_low
+ 7.759000000e-07 V_low
+ 7.759010000e-07 V_hig
+ 7.760000000e-07 V_hig
+ 7.760010000e-07 V_hig
+ 7.761000000e-07 V_hig
+ 7.761010000e-07 V_hig
+ 7.762000000e-07 V_hig
+ 7.762010000e-07 V_hig
+ 7.763000000e-07 V_hig
+ 7.763010000e-07 V_hig
+ 7.764000000e-07 V_hig
+ 7.764010000e-07 V_hig
+ 7.765000000e-07 V_hig
+ 7.765010000e-07 V_hig
+ 7.766000000e-07 V_hig
+ 7.766010000e-07 V_hig
+ 7.767000000e-07 V_hig
+ 7.767010000e-07 V_hig
+ 7.768000000e-07 V_hig
+ 7.768010000e-07 V_hig
+ 7.769000000e-07 V_hig
+ 7.769010000e-07 V_low
+ 7.770000000e-07 V_low
+ 7.770010000e-07 V_low
+ 7.771000000e-07 V_low
+ 7.771010000e-07 V_low
+ 7.772000000e-07 V_low
+ 7.772010000e-07 V_low
+ 7.773000000e-07 V_low
+ 7.773010000e-07 V_low
+ 7.774000000e-07 V_low
+ 7.774010000e-07 V_low
+ 7.775000000e-07 V_low
+ 7.775010000e-07 V_low
+ 7.776000000e-07 V_low
+ 7.776010000e-07 V_low
+ 7.777000000e-07 V_low
+ 7.777010000e-07 V_low
+ 7.778000000e-07 V_low
+ 7.778010000e-07 V_low
+ 7.779000000e-07 V_low
+ 7.779010000e-07 V_low
+ 7.780000000e-07 V_low
+ 7.780010000e-07 V_low
+ 7.781000000e-07 V_low
+ 7.781010000e-07 V_low
+ 7.782000000e-07 V_low
+ 7.782010000e-07 V_low
+ 7.783000000e-07 V_low
+ 7.783010000e-07 V_low
+ 7.784000000e-07 V_low
+ 7.784010000e-07 V_low
+ 7.785000000e-07 V_low
+ 7.785010000e-07 V_low
+ 7.786000000e-07 V_low
+ 7.786010000e-07 V_low
+ 7.787000000e-07 V_low
+ 7.787010000e-07 V_low
+ 7.788000000e-07 V_low
+ 7.788010000e-07 V_low
+ 7.789000000e-07 V_low
+ 7.789010000e-07 V_low
+ 7.790000000e-07 V_low
+ 7.790010000e-07 V_low
+ 7.791000000e-07 V_low
+ 7.791010000e-07 V_low
+ 7.792000000e-07 V_low
+ 7.792010000e-07 V_low
+ 7.793000000e-07 V_low
+ 7.793010000e-07 V_low
+ 7.794000000e-07 V_low
+ 7.794010000e-07 V_low
+ 7.795000000e-07 V_low
+ 7.795010000e-07 V_low
+ 7.796000000e-07 V_low
+ 7.796010000e-07 V_low
+ 7.797000000e-07 V_low
+ 7.797010000e-07 V_low
+ 7.798000000e-07 V_low
+ 7.798010000e-07 V_low
+ 7.799000000e-07 V_low
+ 7.799010000e-07 V_hig
+ 7.800000000e-07 V_hig
+ 7.800010000e-07 V_hig
+ 7.801000000e-07 V_hig
+ 7.801010000e-07 V_hig
+ 7.802000000e-07 V_hig
+ 7.802010000e-07 V_hig
+ 7.803000000e-07 V_hig
+ 7.803010000e-07 V_hig
+ 7.804000000e-07 V_hig
+ 7.804010000e-07 V_hig
+ 7.805000000e-07 V_hig
+ 7.805010000e-07 V_hig
+ 7.806000000e-07 V_hig
+ 7.806010000e-07 V_hig
+ 7.807000000e-07 V_hig
+ 7.807010000e-07 V_hig
+ 7.808000000e-07 V_hig
+ 7.808010000e-07 V_hig
+ 7.809000000e-07 V_hig
+ 7.809010000e-07 V_hig
+ 7.810000000e-07 V_hig
+ 7.810010000e-07 V_hig
+ 7.811000000e-07 V_hig
+ 7.811010000e-07 V_hig
+ 7.812000000e-07 V_hig
+ 7.812010000e-07 V_hig
+ 7.813000000e-07 V_hig
+ 7.813010000e-07 V_hig
+ 7.814000000e-07 V_hig
+ 7.814010000e-07 V_hig
+ 7.815000000e-07 V_hig
+ 7.815010000e-07 V_hig
+ 7.816000000e-07 V_hig
+ 7.816010000e-07 V_hig
+ 7.817000000e-07 V_hig
+ 7.817010000e-07 V_hig
+ 7.818000000e-07 V_hig
+ 7.818010000e-07 V_hig
+ 7.819000000e-07 V_hig
+ 7.819010000e-07 V_hig
+ 7.820000000e-07 V_hig
+ 7.820010000e-07 V_hig
+ 7.821000000e-07 V_hig
+ 7.821010000e-07 V_hig
+ 7.822000000e-07 V_hig
+ 7.822010000e-07 V_hig
+ 7.823000000e-07 V_hig
+ 7.823010000e-07 V_hig
+ 7.824000000e-07 V_hig
+ 7.824010000e-07 V_hig
+ 7.825000000e-07 V_hig
+ 7.825010000e-07 V_hig
+ 7.826000000e-07 V_hig
+ 7.826010000e-07 V_hig
+ 7.827000000e-07 V_hig
+ 7.827010000e-07 V_hig
+ 7.828000000e-07 V_hig
+ 7.828010000e-07 V_hig
+ 7.829000000e-07 V_hig
+ 7.829010000e-07 V_hig
+ 7.830000000e-07 V_hig
+ 7.830010000e-07 V_hig
+ 7.831000000e-07 V_hig
+ 7.831010000e-07 V_hig
+ 7.832000000e-07 V_hig
+ 7.832010000e-07 V_hig
+ 7.833000000e-07 V_hig
+ 7.833010000e-07 V_hig
+ 7.834000000e-07 V_hig
+ 7.834010000e-07 V_hig
+ 7.835000000e-07 V_hig
+ 7.835010000e-07 V_hig
+ 7.836000000e-07 V_hig
+ 7.836010000e-07 V_hig
+ 7.837000000e-07 V_hig
+ 7.837010000e-07 V_hig
+ 7.838000000e-07 V_hig
+ 7.838010000e-07 V_hig
+ 7.839000000e-07 V_hig
+ 7.839010000e-07 V_low
+ 7.840000000e-07 V_low
+ 7.840010000e-07 V_low
+ 7.841000000e-07 V_low
+ 7.841010000e-07 V_low
+ 7.842000000e-07 V_low
+ 7.842010000e-07 V_low
+ 7.843000000e-07 V_low
+ 7.843010000e-07 V_low
+ 7.844000000e-07 V_low
+ 7.844010000e-07 V_low
+ 7.845000000e-07 V_low
+ 7.845010000e-07 V_low
+ 7.846000000e-07 V_low
+ 7.846010000e-07 V_low
+ 7.847000000e-07 V_low
+ 7.847010000e-07 V_low
+ 7.848000000e-07 V_low
+ 7.848010000e-07 V_low
+ 7.849000000e-07 V_low
+ 7.849010000e-07 V_low
+ 7.850000000e-07 V_low
+ 7.850010000e-07 V_low
+ 7.851000000e-07 V_low
+ 7.851010000e-07 V_low
+ 7.852000000e-07 V_low
+ 7.852010000e-07 V_low
+ 7.853000000e-07 V_low
+ 7.853010000e-07 V_low
+ 7.854000000e-07 V_low
+ 7.854010000e-07 V_low
+ 7.855000000e-07 V_low
+ 7.855010000e-07 V_low
+ 7.856000000e-07 V_low
+ 7.856010000e-07 V_low
+ 7.857000000e-07 V_low
+ 7.857010000e-07 V_low
+ 7.858000000e-07 V_low
+ 7.858010000e-07 V_low
+ 7.859000000e-07 V_low
+ 7.859010000e-07 V_hig
+ 7.860000000e-07 V_hig
+ 7.860010000e-07 V_hig
+ 7.861000000e-07 V_hig
+ 7.861010000e-07 V_hig
+ 7.862000000e-07 V_hig
+ 7.862010000e-07 V_hig
+ 7.863000000e-07 V_hig
+ 7.863010000e-07 V_hig
+ 7.864000000e-07 V_hig
+ 7.864010000e-07 V_hig
+ 7.865000000e-07 V_hig
+ 7.865010000e-07 V_hig
+ 7.866000000e-07 V_hig
+ 7.866010000e-07 V_hig
+ 7.867000000e-07 V_hig
+ 7.867010000e-07 V_hig
+ 7.868000000e-07 V_hig
+ 7.868010000e-07 V_hig
+ 7.869000000e-07 V_hig
+ 7.869010000e-07 V_low
+ 7.870000000e-07 V_low
+ 7.870010000e-07 V_low
+ 7.871000000e-07 V_low
+ 7.871010000e-07 V_low
+ 7.872000000e-07 V_low
+ 7.872010000e-07 V_low
+ 7.873000000e-07 V_low
+ 7.873010000e-07 V_low
+ 7.874000000e-07 V_low
+ 7.874010000e-07 V_low
+ 7.875000000e-07 V_low
+ 7.875010000e-07 V_low
+ 7.876000000e-07 V_low
+ 7.876010000e-07 V_low
+ 7.877000000e-07 V_low
+ 7.877010000e-07 V_low
+ 7.878000000e-07 V_low
+ 7.878010000e-07 V_low
+ 7.879000000e-07 V_low
+ 7.879010000e-07 V_hig
+ 7.880000000e-07 V_hig
+ 7.880010000e-07 V_hig
+ 7.881000000e-07 V_hig
+ 7.881010000e-07 V_hig
+ 7.882000000e-07 V_hig
+ 7.882010000e-07 V_hig
+ 7.883000000e-07 V_hig
+ 7.883010000e-07 V_hig
+ 7.884000000e-07 V_hig
+ 7.884010000e-07 V_hig
+ 7.885000000e-07 V_hig
+ 7.885010000e-07 V_hig
+ 7.886000000e-07 V_hig
+ 7.886010000e-07 V_hig
+ 7.887000000e-07 V_hig
+ 7.887010000e-07 V_hig
+ 7.888000000e-07 V_hig
+ 7.888010000e-07 V_hig
+ 7.889000000e-07 V_hig
+ 7.889010000e-07 V_hig
+ 7.890000000e-07 V_hig
+ 7.890010000e-07 V_hig
+ 7.891000000e-07 V_hig
+ 7.891010000e-07 V_hig
+ 7.892000000e-07 V_hig
+ 7.892010000e-07 V_hig
+ 7.893000000e-07 V_hig
+ 7.893010000e-07 V_hig
+ 7.894000000e-07 V_hig
+ 7.894010000e-07 V_hig
+ 7.895000000e-07 V_hig
+ 7.895010000e-07 V_hig
+ 7.896000000e-07 V_hig
+ 7.896010000e-07 V_hig
+ 7.897000000e-07 V_hig
+ 7.897010000e-07 V_hig
+ 7.898000000e-07 V_hig
+ 7.898010000e-07 V_hig
+ 7.899000000e-07 V_hig
+ 7.899010000e-07 V_low
+ 7.900000000e-07 V_low
+ 7.900010000e-07 V_low
+ 7.901000000e-07 V_low
+ 7.901010000e-07 V_low
+ 7.902000000e-07 V_low
+ 7.902010000e-07 V_low
+ 7.903000000e-07 V_low
+ 7.903010000e-07 V_low
+ 7.904000000e-07 V_low
+ 7.904010000e-07 V_low
+ 7.905000000e-07 V_low
+ 7.905010000e-07 V_low
+ 7.906000000e-07 V_low
+ 7.906010000e-07 V_low
+ 7.907000000e-07 V_low
+ 7.907010000e-07 V_low
+ 7.908000000e-07 V_low
+ 7.908010000e-07 V_low
+ 7.909000000e-07 V_low
+ 7.909010000e-07 V_low
+ 7.910000000e-07 V_low
+ 7.910010000e-07 V_low
+ 7.911000000e-07 V_low
+ 7.911010000e-07 V_low
+ 7.912000000e-07 V_low
+ 7.912010000e-07 V_low
+ 7.913000000e-07 V_low
+ 7.913010000e-07 V_low
+ 7.914000000e-07 V_low
+ 7.914010000e-07 V_low
+ 7.915000000e-07 V_low
+ 7.915010000e-07 V_low
+ 7.916000000e-07 V_low
+ 7.916010000e-07 V_low
+ 7.917000000e-07 V_low
+ 7.917010000e-07 V_low
+ 7.918000000e-07 V_low
+ 7.918010000e-07 V_low
+ 7.919000000e-07 V_low
+ 7.919010000e-07 V_low
+ 7.920000000e-07 V_low
+ 7.920010000e-07 V_low
+ 7.921000000e-07 V_low
+ 7.921010000e-07 V_low
+ 7.922000000e-07 V_low
+ 7.922010000e-07 V_low
+ 7.923000000e-07 V_low
+ 7.923010000e-07 V_low
+ 7.924000000e-07 V_low
+ 7.924010000e-07 V_low
+ 7.925000000e-07 V_low
+ 7.925010000e-07 V_low
+ 7.926000000e-07 V_low
+ 7.926010000e-07 V_low
+ 7.927000000e-07 V_low
+ 7.927010000e-07 V_low
+ 7.928000000e-07 V_low
+ 7.928010000e-07 V_low
+ 7.929000000e-07 V_low
+ 7.929010000e-07 V_low
+ 7.930000000e-07 V_low
+ 7.930010000e-07 V_low
+ 7.931000000e-07 V_low
+ 7.931010000e-07 V_low
+ 7.932000000e-07 V_low
+ 7.932010000e-07 V_low
+ 7.933000000e-07 V_low
+ 7.933010000e-07 V_low
+ 7.934000000e-07 V_low
+ 7.934010000e-07 V_low
+ 7.935000000e-07 V_low
+ 7.935010000e-07 V_low
+ 7.936000000e-07 V_low
+ 7.936010000e-07 V_low
+ 7.937000000e-07 V_low
+ 7.937010000e-07 V_low
+ 7.938000000e-07 V_low
+ 7.938010000e-07 V_low
+ 7.939000000e-07 V_low
+ 7.939010000e-07 V_low
+ 7.940000000e-07 V_low
+ 7.940010000e-07 V_low
+ 7.941000000e-07 V_low
+ 7.941010000e-07 V_low
+ 7.942000000e-07 V_low
+ 7.942010000e-07 V_low
+ 7.943000000e-07 V_low
+ 7.943010000e-07 V_low
+ 7.944000000e-07 V_low
+ 7.944010000e-07 V_low
+ 7.945000000e-07 V_low
+ 7.945010000e-07 V_low
+ 7.946000000e-07 V_low
+ 7.946010000e-07 V_low
+ 7.947000000e-07 V_low
+ 7.947010000e-07 V_low
+ 7.948000000e-07 V_low
+ 7.948010000e-07 V_low
+ 7.949000000e-07 V_low
+ 7.949010000e-07 V_hig
+ 7.950000000e-07 V_hig
+ 7.950010000e-07 V_hig
+ 7.951000000e-07 V_hig
+ 7.951010000e-07 V_hig
+ 7.952000000e-07 V_hig
+ 7.952010000e-07 V_hig
+ 7.953000000e-07 V_hig
+ 7.953010000e-07 V_hig
+ 7.954000000e-07 V_hig
+ 7.954010000e-07 V_hig
+ 7.955000000e-07 V_hig
+ 7.955010000e-07 V_hig
+ 7.956000000e-07 V_hig
+ 7.956010000e-07 V_hig
+ 7.957000000e-07 V_hig
+ 7.957010000e-07 V_hig
+ 7.958000000e-07 V_hig
+ 7.958010000e-07 V_hig
+ 7.959000000e-07 V_hig
+ 7.959010000e-07 V_low
+ 7.960000000e-07 V_low
+ 7.960010000e-07 V_low
+ 7.961000000e-07 V_low
+ 7.961010000e-07 V_low
+ 7.962000000e-07 V_low
+ 7.962010000e-07 V_low
+ 7.963000000e-07 V_low
+ 7.963010000e-07 V_low
+ 7.964000000e-07 V_low
+ 7.964010000e-07 V_low
+ 7.965000000e-07 V_low
+ 7.965010000e-07 V_low
+ 7.966000000e-07 V_low
+ 7.966010000e-07 V_low
+ 7.967000000e-07 V_low
+ 7.967010000e-07 V_low
+ 7.968000000e-07 V_low
+ 7.968010000e-07 V_low
+ 7.969000000e-07 V_low
+ 7.969010000e-07 V_hig
+ 7.970000000e-07 V_hig
+ 7.970010000e-07 V_hig
+ 7.971000000e-07 V_hig
+ 7.971010000e-07 V_hig
+ 7.972000000e-07 V_hig
+ 7.972010000e-07 V_hig
+ 7.973000000e-07 V_hig
+ 7.973010000e-07 V_hig
+ 7.974000000e-07 V_hig
+ 7.974010000e-07 V_hig
+ 7.975000000e-07 V_hig
+ 7.975010000e-07 V_hig
+ 7.976000000e-07 V_hig
+ 7.976010000e-07 V_hig
+ 7.977000000e-07 V_hig
+ 7.977010000e-07 V_hig
+ 7.978000000e-07 V_hig
+ 7.978010000e-07 V_hig
+ 7.979000000e-07 V_hig
+ 7.979010000e-07 V_low
+ 7.980000000e-07 V_low
+ 7.980010000e-07 V_low
+ 7.981000000e-07 V_low
+ 7.981010000e-07 V_low
+ 7.982000000e-07 V_low
+ 7.982010000e-07 V_low
+ 7.983000000e-07 V_low
+ 7.983010000e-07 V_low
+ 7.984000000e-07 V_low
+ 7.984010000e-07 V_low
+ 7.985000000e-07 V_low
+ 7.985010000e-07 V_low
+ 7.986000000e-07 V_low
+ 7.986010000e-07 V_low
+ 7.987000000e-07 V_low
+ 7.987010000e-07 V_low
+ 7.988000000e-07 V_low
+ 7.988010000e-07 V_low
+ 7.989000000e-07 V_low
+ 7.989010000e-07 V_hig
+ 7.990000000e-07 V_hig
+ 7.990010000e-07 V_hig
+ 7.991000000e-07 V_hig
+ 7.991010000e-07 V_hig
+ 7.992000000e-07 V_hig
+ 7.992010000e-07 V_hig
+ 7.993000000e-07 V_hig
+ 7.993010000e-07 V_hig
+ 7.994000000e-07 V_hig
+ 7.994010000e-07 V_hig
+ 7.995000000e-07 V_hig
+ 7.995010000e-07 V_hig
+ 7.996000000e-07 V_hig
+ 7.996010000e-07 V_hig
+ 7.997000000e-07 V_hig
+ 7.997010000e-07 V_hig
+ 7.998000000e-07 V_hig
+ 7.998010000e-07 V_hig
+ 7.999000000e-07 V_hig
+ 7.999010000e-07 V_hig
+ 8.000000000e-07 V_hig
+ 8.000010000e-07 V_hig
+ 8.001000000e-07 V_hig
+ 8.001010000e-07 V_hig
+ 8.002000000e-07 V_hig
+ 8.002010000e-07 V_hig
+ 8.003000000e-07 V_hig
+ 8.003010000e-07 V_hig
+ 8.004000000e-07 V_hig
+ 8.004010000e-07 V_hig
+ 8.005000000e-07 V_hig
+ 8.005010000e-07 V_hig
+ 8.006000000e-07 V_hig
+ 8.006010000e-07 V_hig
+ 8.007000000e-07 V_hig
+ 8.007010000e-07 V_hig
+ 8.008000000e-07 V_hig
+ 8.008010000e-07 V_hig
+ 8.009000000e-07 V_hig
+ 8.009010000e-07 V_low
+ 8.010000000e-07 V_low
+ 8.010010000e-07 V_low
+ 8.011000000e-07 V_low
+ 8.011010000e-07 V_low
+ 8.012000000e-07 V_low
+ 8.012010000e-07 V_low
+ 8.013000000e-07 V_low
+ 8.013010000e-07 V_low
+ 8.014000000e-07 V_low
+ 8.014010000e-07 V_low
+ 8.015000000e-07 V_low
+ 8.015010000e-07 V_low
+ 8.016000000e-07 V_low
+ 8.016010000e-07 V_low
+ 8.017000000e-07 V_low
+ 8.017010000e-07 V_low
+ 8.018000000e-07 V_low
+ 8.018010000e-07 V_low
+ 8.019000000e-07 V_low
+ 8.019010000e-07 V_low
+ 8.020000000e-07 V_low
+ 8.020010000e-07 V_low
+ 8.021000000e-07 V_low
+ 8.021010000e-07 V_low
+ 8.022000000e-07 V_low
+ 8.022010000e-07 V_low
+ 8.023000000e-07 V_low
+ 8.023010000e-07 V_low
+ 8.024000000e-07 V_low
+ 8.024010000e-07 V_low
+ 8.025000000e-07 V_low
+ 8.025010000e-07 V_low
+ 8.026000000e-07 V_low
+ 8.026010000e-07 V_low
+ 8.027000000e-07 V_low
+ 8.027010000e-07 V_low
+ 8.028000000e-07 V_low
+ 8.028010000e-07 V_low
+ 8.029000000e-07 V_low
+ 8.029010000e-07 V_hig
+ 8.030000000e-07 V_hig
+ 8.030010000e-07 V_hig
+ 8.031000000e-07 V_hig
+ 8.031010000e-07 V_hig
+ 8.032000000e-07 V_hig
+ 8.032010000e-07 V_hig
+ 8.033000000e-07 V_hig
+ 8.033010000e-07 V_hig
+ 8.034000000e-07 V_hig
+ 8.034010000e-07 V_hig
+ 8.035000000e-07 V_hig
+ 8.035010000e-07 V_hig
+ 8.036000000e-07 V_hig
+ 8.036010000e-07 V_hig
+ 8.037000000e-07 V_hig
+ 8.037010000e-07 V_hig
+ 8.038000000e-07 V_hig
+ 8.038010000e-07 V_hig
+ 8.039000000e-07 V_hig
+ 8.039010000e-07 V_low
+ 8.040000000e-07 V_low
+ 8.040010000e-07 V_low
+ 8.041000000e-07 V_low
+ 8.041010000e-07 V_low
+ 8.042000000e-07 V_low
+ 8.042010000e-07 V_low
+ 8.043000000e-07 V_low
+ 8.043010000e-07 V_low
+ 8.044000000e-07 V_low
+ 8.044010000e-07 V_low
+ 8.045000000e-07 V_low
+ 8.045010000e-07 V_low
+ 8.046000000e-07 V_low
+ 8.046010000e-07 V_low
+ 8.047000000e-07 V_low
+ 8.047010000e-07 V_low
+ 8.048000000e-07 V_low
+ 8.048010000e-07 V_low
+ 8.049000000e-07 V_low
+ 8.049010000e-07 V_low
+ 8.050000000e-07 V_low
+ 8.050010000e-07 V_low
+ 8.051000000e-07 V_low
+ 8.051010000e-07 V_low
+ 8.052000000e-07 V_low
+ 8.052010000e-07 V_low
+ 8.053000000e-07 V_low
+ 8.053010000e-07 V_low
+ 8.054000000e-07 V_low
+ 8.054010000e-07 V_low
+ 8.055000000e-07 V_low
+ 8.055010000e-07 V_low
+ 8.056000000e-07 V_low
+ 8.056010000e-07 V_low
+ 8.057000000e-07 V_low
+ 8.057010000e-07 V_low
+ 8.058000000e-07 V_low
+ 8.058010000e-07 V_low
+ 8.059000000e-07 V_low
+ 8.059010000e-07 V_hig
+ 8.060000000e-07 V_hig
+ 8.060010000e-07 V_hig
+ 8.061000000e-07 V_hig
+ 8.061010000e-07 V_hig
+ 8.062000000e-07 V_hig
+ 8.062010000e-07 V_hig
+ 8.063000000e-07 V_hig
+ 8.063010000e-07 V_hig
+ 8.064000000e-07 V_hig
+ 8.064010000e-07 V_hig
+ 8.065000000e-07 V_hig
+ 8.065010000e-07 V_hig
+ 8.066000000e-07 V_hig
+ 8.066010000e-07 V_hig
+ 8.067000000e-07 V_hig
+ 8.067010000e-07 V_hig
+ 8.068000000e-07 V_hig
+ 8.068010000e-07 V_hig
+ 8.069000000e-07 V_hig
+ 8.069010000e-07 V_low
+ 8.070000000e-07 V_low
+ 8.070010000e-07 V_low
+ 8.071000000e-07 V_low
+ 8.071010000e-07 V_low
+ 8.072000000e-07 V_low
+ 8.072010000e-07 V_low
+ 8.073000000e-07 V_low
+ 8.073010000e-07 V_low
+ 8.074000000e-07 V_low
+ 8.074010000e-07 V_low
+ 8.075000000e-07 V_low
+ 8.075010000e-07 V_low
+ 8.076000000e-07 V_low
+ 8.076010000e-07 V_low
+ 8.077000000e-07 V_low
+ 8.077010000e-07 V_low
+ 8.078000000e-07 V_low
+ 8.078010000e-07 V_low
+ 8.079000000e-07 V_low
+ 8.079010000e-07 V_hig
+ 8.080000000e-07 V_hig
+ 8.080010000e-07 V_hig
+ 8.081000000e-07 V_hig
+ 8.081010000e-07 V_hig
+ 8.082000000e-07 V_hig
+ 8.082010000e-07 V_hig
+ 8.083000000e-07 V_hig
+ 8.083010000e-07 V_hig
+ 8.084000000e-07 V_hig
+ 8.084010000e-07 V_hig
+ 8.085000000e-07 V_hig
+ 8.085010000e-07 V_hig
+ 8.086000000e-07 V_hig
+ 8.086010000e-07 V_hig
+ 8.087000000e-07 V_hig
+ 8.087010000e-07 V_hig
+ 8.088000000e-07 V_hig
+ 8.088010000e-07 V_hig
+ 8.089000000e-07 V_hig
+ 8.089010000e-07 V_low
+ 8.090000000e-07 V_low
+ 8.090010000e-07 V_low
+ 8.091000000e-07 V_low
+ 8.091010000e-07 V_low
+ 8.092000000e-07 V_low
+ 8.092010000e-07 V_low
+ 8.093000000e-07 V_low
+ 8.093010000e-07 V_low
+ 8.094000000e-07 V_low
+ 8.094010000e-07 V_low
+ 8.095000000e-07 V_low
+ 8.095010000e-07 V_low
+ 8.096000000e-07 V_low
+ 8.096010000e-07 V_low
+ 8.097000000e-07 V_low
+ 8.097010000e-07 V_low
+ 8.098000000e-07 V_low
+ 8.098010000e-07 V_low
+ 8.099000000e-07 V_low
+ 8.099010000e-07 V_hig
+ 8.100000000e-07 V_hig
+ 8.100010000e-07 V_hig
+ 8.101000000e-07 V_hig
+ 8.101010000e-07 V_hig
+ 8.102000000e-07 V_hig
+ 8.102010000e-07 V_hig
+ 8.103000000e-07 V_hig
+ 8.103010000e-07 V_hig
+ 8.104000000e-07 V_hig
+ 8.104010000e-07 V_hig
+ 8.105000000e-07 V_hig
+ 8.105010000e-07 V_hig
+ 8.106000000e-07 V_hig
+ 8.106010000e-07 V_hig
+ 8.107000000e-07 V_hig
+ 8.107010000e-07 V_hig
+ 8.108000000e-07 V_hig
+ 8.108010000e-07 V_hig
+ 8.109000000e-07 V_hig
+ 8.109010000e-07 V_low
+ 8.110000000e-07 V_low
+ 8.110010000e-07 V_low
+ 8.111000000e-07 V_low
+ 8.111010000e-07 V_low
+ 8.112000000e-07 V_low
+ 8.112010000e-07 V_low
+ 8.113000000e-07 V_low
+ 8.113010000e-07 V_low
+ 8.114000000e-07 V_low
+ 8.114010000e-07 V_low
+ 8.115000000e-07 V_low
+ 8.115010000e-07 V_low
+ 8.116000000e-07 V_low
+ 8.116010000e-07 V_low
+ 8.117000000e-07 V_low
+ 8.117010000e-07 V_low
+ 8.118000000e-07 V_low
+ 8.118010000e-07 V_low
+ 8.119000000e-07 V_low
+ 8.119010000e-07 V_low
+ 8.120000000e-07 V_low
+ 8.120010000e-07 V_low
+ 8.121000000e-07 V_low
+ 8.121010000e-07 V_low
+ 8.122000000e-07 V_low
+ 8.122010000e-07 V_low
+ 8.123000000e-07 V_low
+ 8.123010000e-07 V_low
+ 8.124000000e-07 V_low
+ 8.124010000e-07 V_low
+ 8.125000000e-07 V_low
+ 8.125010000e-07 V_low
+ 8.126000000e-07 V_low
+ 8.126010000e-07 V_low
+ 8.127000000e-07 V_low
+ 8.127010000e-07 V_low
+ 8.128000000e-07 V_low
+ 8.128010000e-07 V_low
+ 8.129000000e-07 V_low
+ 8.129010000e-07 V_low
+ 8.130000000e-07 V_low
+ 8.130010000e-07 V_low
+ 8.131000000e-07 V_low
+ 8.131010000e-07 V_low
+ 8.132000000e-07 V_low
+ 8.132010000e-07 V_low
+ 8.133000000e-07 V_low
+ 8.133010000e-07 V_low
+ 8.134000000e-07 V_low
+ 8.134010000e-07 V_low
+ 8.135000000e-07 V_low
+ 8.135010000e-07 V_low
+ 8.136000000e-07 V_low
+ 8.136010000e-07 V_low
+ 8.137000000e-07 V_low
+ 8.137010000e-07 V_low
+ 8.138000000e-07 V_low
+ 8.138010000e-07 V_low
+ 8.139000000e-07 V_low
+ 8.139010000e-07 V_hig
+ 8.140000000e-07 V_hig
+ 8.140010000e-07 V_hig
+ 8.141000000e-07 V_hig
+ 8.141010000e-07 V_hig
+ 8.142000000e-07 V_hig
+ 8.142010000e-07 V_hig
+ 8.143000000e-07 V_hig
+ 8.143010000e-07 V_hig
+ 8.144000000e-07 V_hig
+ 8.144010000e-07 V_hig
+ 8.145000000e-07 V_hig
+ 8.145010000e-07 V_hig
+ 8.146000000e-07 V_hig
+ 8.146010000e-07 V_hig
+ 8.147000000e-07 V_hig
+ 8.147010000e-07 V_hig
+ 8.148000000e-07 V_hig
+ 8.148010000e-07 V_hig
+ 8.149000000e-07 V_hig
+ 8.149010000e-07 V_low
+ 8.150000000e-07 V_low
+ 8.150010000e-07 V_low
+ 8.151000000e-07 V_low
+ 8.151010000e-07 V_low
+ 8.152000000e-07 V_low
+ 8.152010000e-07 V_low
+ 8.153000000e-07 V_low
+ 8.153010000e-07 V_low
+ 8.154000000e-07 V_low
+ 8.154010000e-07 V_low
+ 8.155000000e-07 V_low
+ 8.155010000e-07 V_low
+ 8.156000000e-07 V_low
+ 8.156010000e-07 V_low
+ 8.157000000e-07 V_low
+ 8.157010000e-07 V_low
+ 8.158000000e-07 V_low
+ 8.158010000e-07 V_low
+ 8.159000000e-07 V_low
+ 8.159010000e-07 V_hig
+ 8.160000000e-07 V_hig
+ 8.160010000e-07 V_hig
+ 8.161000000e-07 V_hig
+ 8.161010000e-07 V_hig
+ 8.162000000e-07 V_hig
+ 8.162010000e-07 V_hig
+ 8.163000000e-07 V_hig
+ 8.163010000e-07 V_hig
+ 8.164000000e-07 V_hig
+ 8.164010000e-07 V_hig
+ 8.165000000e-07 V_hig
+ 8.165010000e-07 V_hig
+ 8.166000000e-07 V_hig
+ 8.166010000e-07 V_hig
+ 8.167000000e-07 V_hig
+ 8.167010000e-07 V_hig
+ 8.168000000e-07 V_hig
+ 8.168010000e-07 V_hig
+ 8.169000000e-07 V_hig
+ 8.169010000e-07 V_low
+ 8.170000000e-07 V_low
+ 8.170010000e-07 V_low
+ 8.171000000e-07 V_low
+ 8.171010000e-07 V_low
+ 8.172000000e-07 V_low
+ 8.172010000e-07 V_low
+ 8.173000000e-07 V_low
+ 8.173010000e-07 V_low
+ 8.174000000e-07 V_low
+ 8.174010000e-07 V_low
+ 8.175000000e-07 V_low
+ 8.175010000e-07 V_low
+ 8.176000000e-07 V_low
+ 8.176010000e-07 V_low
+ 8.177000000e-07 V_low
+ 8.177010000e-07 V_low
+ 8.178000000e-07 V_low
+ 8.178010000e-07 V_low
+ 8.179000000e-07 V_low
+ 8.179010000e-07 V_low
+ 8.180000000e-07 V_low
+ 8.180010000e-07 V_low
+ 8.181000000e-07 V_low
+ 8.181010000e-07 V_low
+ 8.182000000e-07 V_low
+ 8.182010000e-07 V_low
+ 8.183000000e-07 V_low
+ 8.183010000e-07 V_low
+ 8.184000000e-07 V_low
+ 8.184010000e-07 V_low
+ 8.185000000e-07 V_low
+ 8.185010000e-07 V_low
+ 8.186000000e-07 V_low
+ 8.186010000e-07 V_low
+ 8.187000000e-07 V_low
+ 8.187010000e-07 V_low
+ 8.188000000e-07 V_low
+ 8.188010000e-07 V_low
+ 8.189000000e-07 V_low
+ 8.189010000e-07 V_hig
+ 8.190000000e-07 V_hig
+ 8.190010000e-07 V_hig
+ 8.191000000e-07 V_hig
+ 8.191010000e-07 V_hig
+ 8.192000000e-07 V_hig
+ 8.192010000e-07 V_hig
+ 8.193000000e-07 V_hig
+ 8.193010000e-07 V_hig
+ 8.194000000e-07 V_hig
+ 8.194010000e-07 V_hig
+ 8.195000000e-07 V_hig
+ 8.195010000e-07 V_hig
+ 8.196000000e-07 V_hig
+ 8.196010000e-07 V_hig
+ 8.197000000e-07 V_hig
+ 8.197010000e-07 V_hig
+ 8.198000000e-07 V_hig
+ 8.198010000e-07 V_hig
+ 8.199000000e-07 V_hig
+ 8.199010000e-07 V_low
+ 8.200000000e-07 V_low
+ 8.200010000e-07 V_low
+ 8.201000000e-07 V_low
+ 8.201010000e-07 V_low
+ 8.202000000e-07 V_low
+ 8.202010000e-07 V_low
+ 8.203000000e-07 V_low
+ 8.203010000e-07 V_low
+ 8.204000000e-07 V_low
+ 8.204010000e-07 V_low
+ 8.205000000e-07 V_low
+ 8.205010000e-07 V_low
+ 8.206000000e-07 V_low
+ 8.206010000e-07 V_low
+ 8.207000000e-07 V_low
+ 8.207010000e-07 V_low
+ 8.208000000e-07 V_low
+ 8.208010000e-07 V_low
+ 8.209000000e-07 V_low
+ 8.209010000e-07 V_low
+ 8.210000000e-07 V_low
+ 8.210010000e-07 V_low
+ 8.211000000e-07 V_low
+ 8.211010000e-07 V_low
+ 8.212000000e-07 V_low
+ 8.212010000e-07 V_low
+ 8.213000000e-07 V_low
+ 8.213010000e-07 V_low
+ 8.214000000e-07 V_low
+ 8.214010000e-07 V_low
+ 8.215000000e-07 V_low
+ 8.215010000e-07 V_low
+ 8.216000000e-07 V_low
+ 8.216010000e-07 V_low
+ 8.217000000e-07 V_low
+ 8.217010000e-07 V_low
+ 8.218000000e-07 V_low
+ 8.218010000e-07 V_low
+ 8.219000000e-07 V_low
+ 8.219010000e-07 V_low
+ 8.220000000e-07 V_low
+ 8.220010000e-07 V_low
+ 8.221000000e-07 V_low
+ 8.221010000e-07 V_low
+ 8.222000000e-07 V_low
+ 8.222010000e-07 V_low
+ 8.223000000e-07 V_low
+ 8.223010000e-07 V_low
+ 8.224000000e-07 V_low
+ 8.224010000e-07 V_low
+ 8.225000000e-07 V_low
+ 8.225010000e-07 V_low
+ 8.226000000e-07 V_low
+ 8.226010000e-07 V_low
+ 8.227000000e-07 V_low
+ 8.227010000e-07 V_low
+ 8.228000000e-07 V_low
+ 8.228010000e-07 V_low
+ 8.229000000e-07 V_low
+ 8.229010000e-07 V_hig
+ 8.230000000e-07 V_hig
+ 8.230010000e-07 V_hig
+ 8.231000000e-07 V_hig
+ 8.231010000e-07 V_hig
+ 8.232000000e-07 V_hig
+ 8.232010000e-07 V_hig
+ 8.233000000e-07 V_hig
+ 8.233010000e-07 V_hig
+ 8.234000000e-07 V_hig
+ 8.234010000e-07 V_hig
+ 8.235000000e-07 V_hig
+ 8.235010000e-07 V_hig
+ 8.236000000e-07 V_hig
+ 8.236010000e-07 V_hig
+ 8.237000000e-07 V_hig
+ 8.237010000e-07 V_hig
+ 8.238000000e-07 V_hig
+ 8.238010000e-07 V_hig
+ 8.239000000e-07 V_hig
+ 8.239010000e-07 V_low
+ 8.240000000e-07 V_low
+ 8.240010000e-07 V_low
+ 8.241000000e-07 V_low
+ 8.241010000e-07 V_low
+ 8.242000000e-07 V_low
+ 8.242010000e-07 V_low
+ 8.243000000e-07 V_low
+ 8.243010000e-07 V_low
+ 8.244000000e-07 V_low
+ 8.244010000e-07 V_low
+ 8.245000000e-07 V_low
+ 8.245010000e-07 V_low
+ 8.246000000e-07 V_low
+ 8.246010000e-07 V_low
+ 8.247000000e-07 V_low
+ 8.247010000e-07 V_low
+ 8.248000000e-07 V_low
+ 8.248010000e-07 V_low
+ 8.249000000e-07 V_low
+ 8.249010000e-07 V_low
+ 8.250000000e-07 V_low
+ 8.250010000e-07 V_low
+ 8.251000000e-07 V_low
+ 8.251010000e-07 V_low
+ 8.252000000e-07 V_low
+ 8.252010000e-07 V_low
+ 8.253000000e-07 V_low
+ 8.253010000e-07 V_low
+ 8.254000000e-07 V_low
+ 8.254010000e-07 V_low
+ 8.255000000e-07 V_low
+ 8.255010000e-07 V_low
+ 8.256000000e-07 V_low
+ 8.256010000e-07 V_low
+ 8.257000000e-07 V_low
+ 8.257010000e-07 V_low
+ 8.258000000e-07 V_low
+ 8.258010000e-07 V_low
+ 8.259000000e-07 V_low
+ 8.259010000e-07 V_hig
+ 8.260000000e-07 V_hig
+ 8.260010000e-07 V_hig
+ 8.261000000e-07 V_hig
+ 8.261010000e-07 V_hig
+ 8.262000000e-07 V_hig
+ 8.262010000e-07 V_hig
+ 8.263000000e-07 V_hig
+ 8.263010000e-07 V_hig
+ 8.264000000e-07 V_hig
+ 8.264010000e-07 V_hig
+ 8.265000000e-07 V_hig
+ 8.265010000e-07 V_hig
+ 8.266000000e-07 V_hig
+ 8.266010000e-07 V_hig
+ 8.267000000e-07 V_hig
+ 8.267010000e-07 V_hig
+ 8.268000000e-07 V_hig
+ 8.268010000e-07 V_hig
+ 8.269000000e-07 V_hig
+ 8.269010000e-07 V_hig
+ 8.270000000e-07 V_hig
+ 8.270010000e-07 V_hig
+ 8.271000000e-07 V_hig
+ 8.271010000e-07 V_hig
+ 8.272000000e-07 V_hig
+ 8.272010000e-07 V_hig
+ 8.273000000e-07 V_hig
+ 8.273010000e-07 V_hig
+ 8.274000000e-07 V_hig
+ 8.274010000e-07 V_hig
+ 8.275000000e-07 V_hig
+ 8.275010000e-07 V_hig
+ 8.276000000e-07 V_hig
+ 8.276010000e-07 V_hig
+ 8.277000000e-07 V_hig
+ 8.277010000e-07 V_hig
+ 8.278000000e-07 V_hig
+ 8.278010000e-07 V_hig
+ 8.279000000e-07 V_hig
+ 8.279010000e-07 V_low
+ 8.280000000e-07 V_low
+ 8.280010000e-07 V_low
+ 8.281000000e-07 V_low
+ 8.281010000e-07 V_low
+ 8.282000000e-07 V_low
+ 8.282010000e-07 V_low
+ 8.283000000e-07 V_low
+ 8.283010000e-07 V_low
+ 8.284000000e-07 V_low
+ 8.284010000e-07 V_low
+ 8.285000000e-07 V_low
+ 8.285010000e-07 V_low
+ 8.286000000e-07 V_low
+ 8.286010000e-07 V_low
+ 8.287000000e-07 V_low
+ 8.287010000e-07 V_low
+ 8.288000000e-07 V_low
+ 8.288010000e-07 V_low
+ 8.289000000e-07 V_low
+ 8.289010000e-07 V_hig
+ 8.290000000e-07 V_hig
+ 8.290010000e-07 V_hig
+ 8.291000000e-07 V_hig
+ 8.291010000e-07 V_hig
+ 8.292000000e-07 V_hig
+ 8.292010000e-07 V_hig
+ 8.293000000e-07 V_hig
+ 8.293010000e-07 V_hig
+ 8.294000000e-07 V_hig
+ 8.294010000e-07 V_hig
+ 8.295000000e-07 V_hig
+ 8.295010000e-07 V_hig
+ 8.296000000e-07 V_hig
+ 8.296010000e-07 V_hig
+ 8.297000000e-07 V_hig
+ 8.297010000e-07 V_hig
+ 8.298000000e-07 V_hig
+ 8.298010000e-07 V_hig
+ 8.299000000e-07 V_hig
+ 8.299010000e-07 V_hig
+ 8.300000000e-07 V_hig
+ 8.300010000e-07 V_hig
+ 8.301000000e-07 V_hig
+ 8.301010000e-07 V_hig
+ 8.302000000e-07 V_hig
+ 8.302010000e-07 V_hig
+ 8.303000000e-07 V_hig
+ 8.303010000e-07 V_hig
+ 8.304000000e-07 V_hig
+ 8.304010000e-07 V_hig
+ 8.305000000e-07 V_hig
+ 8.305010000e-07 V_hig
+ 8.306000000e-07 V_hig
+ 8.306010000e-07 V_hig
+ 8.307000000e-07 V_hig
+ 8.307010000e-07 V_hig
+ 8.308000000e-07 V_hig
+ 8.308010000e-07 V_hig
+ 8.309000000e-07 V_hig
+ 8.309010000e-07 V_hig
+ 8.310000000e-07 V_hig
+ 8.310010000e-07 V_hig
+ 8.311000000e-07 V_hig
+ 8.311010000e-07 V_hig
+ 8.312000000e-07 V_hig
+ 8.312010000e-07 V_hig
+ 8.313000000e-07 V_hig
+ 8.313010000e-07 V_hig
+ 8.314000000e-07 V_hig
+ 8.314010000e-07 V_hig
+ 8.315000000e-07 V_hig
+ 8.315010000e-07 V_hig
+ 8.316000000e-07 V_hig
+ 8.316010000e-07 V_hig
+ 8.317000000e-07 V_hig
+ 8.317010000e-07 V_hig
+ 8.318000000e-07 V_hig
+ 8.318010000e-07 V_hig
+ 8.319000000e-07 V_hig
+ 8.319010000e-07 V_low
+ 8.320000000e-07 V_low
+ 8.320010000e-07 V_low
+ 8.321000000e-07 V_low
+ 8.321010000e-07 V_low
+ 8.322000000e-07 V_low
+ 8.322010000e-07 V_low
+ 8.323000000e-07 V_low
+ 8.323010000e-07 V_low
+ 8.324000000e-07 V_low
+ 8.324010000e-07 V_low
+ 8.325000000e-07 V_low
+ 8.325010000e-07 V_low
+ 8.326000000e-07 V_low
+ 8.326010000e-07 V_low
+ 8.327000000e-07 V_low
+ 8.327010000e-07 V_low
+ 8.328000000e-07 V_low
+ 8.328010000e-07 V_low
+ 8.329000000e-07 V_low
+ 8.329010000e-07 V_low
+ 8.330000000e-07 V_low
+ 8.330010000e-07 V_low
+ 8.331000000e-07 V_low
+ 8.331010000e-07 V_low
+ 8.332000000e-07 V_low
+ 8.332010000e-07 V_low
+ 8.333000000e-07 V_low
+ 8.333010000e-07 V_low
+ 8.334000000e-07 V_low
+ 8.334010000e-07 V_low
+ 8.335000000e-07 V_low
+ 8.335010000e-07 V_low
+ 8.336000000e-07 V_low
+ 8.336010000e-07 V_low
+ 8.337000000e-07 V_low
+ 8.337010000e-07 V_low
+ 8.338000000e-07 V_low
+ 8.338010000e-07 V_low
+ 8.339000000e-07 V_low
+ 8.339010000e-07 V_hig
+ 8.340000000e-07 V_hig
+ 8.340010000e-07 V_hig
+ 8.341000000e-07 V_hig
+ 8.341010000e-07 V_hig
+ 8.342000000e-07 V_hig
+ 8.342010000e-07 V_hig
+ 8.343000000e-07 V_hig
+ 8.343010000e-07 V_hig
+ 8.344000000e-07 V_hig
+ 8.344010000e-07 V_hig
+ 8.345000000e-07 V_hig
+ 8.345010000e-07 V_hig
+ 8.346000000e-07 V_hig
+ 8.346010000e-07 V_hig
+ 8.347000000e-07 V_hig
+ 8.347010000e-07 V_hig
+ 8.348000000e-07 V_hig
+ 8.348010000e-07 V_hig
+ 8.349000000e-07 V_hig
+ 8.349010000e-07 V_hig
+ 8.350000000e-07 V_hig
+ 8.350010000e-07 V_hig
+ 8.351000000e-07 V_hig
+ 8.351010000e-07 V_hig
+ 8.352000000e-07 V_hig
+ 8.352010000e-07 V_hig
+ 8.353000000e-07 V_hig
+ 8.353010000e-07 V_hig
+ 8.354000000e-07 V_hig
+ 8.354010000e-07 V_hig
+ 8.355000000e-07 V_hig
+ 8.355010000e-07 V_hig
+ 8.356000000e-07 V_hig
+ 8.356010000e-07 V_hig
+ 8.357000000e-07 V_hig
+ 8.357010000e-07 V_hig
+ 8.358000000e-07 V_hig
+ 8.358010000e-07 V_hig
+ 8.359000000e-07 V_hig
+ 8.359010000e-07 V_low
+ 8.360000000e-07 V_low
+ 8.360010000e-07 V_low
+ 8.361000000e-07 V_low
+ 8.361010000e-07 V_low
+ 8.362000000e-07 V_low
+ 8.362010000e-07 V_low
+ 8.363000000e-07 V_low
+ 8.363010000e-07 V_low
+ 8.364000000e-07 V_low
+ 8.364010000e-07 V_low
+ 8.365000000e-07 V_low
+ 8.365010000e-07 V_low
+ 8.366000000e-07 V_low
+ 8.366010000e-07 V_low
+ 8.367000000e-07 V_low
+ 8.367010000e-07 V_low
+ 8.368000000e-07 V_low
+ 8.368010000e-07 V_low
+ 8.369000000e-07 V_low
+ 8.369010000e-07 V_low
+ 8.370000000e-07 V_low
+ 8.370010000e-07 V_low
+ 8.371000000e-07 V_low
+ 8.371010000e-07 V_low
+ 8.372000000e-07 V_low
+ 8.372010000e-07 V_low
+ 8.373000000e-07 V_low
+ 8.373010000e-07 V_low
+ 8.374000000e-07 V_low
+ 8.374010000e-07 V_low
+ 8.375000000e-07 V_low
+ 8.375010000e-07 V_low
+ 8.376000000e-07 V_low
+ 8.376010000e-07 V_low
+ 8.377000000e-07 V_low
+ 8.377010000e-07 V_low
+ 8.378000000e-07 V_low
+ 8.378010000e-07 V_low
+ 8.379000000e-07 V_low
+ 8.379010000e-07 V_low
+ 8.380000000e-07 V_low
+ 8.380010000e-07 V_low
+ 8.381000000e-07 V_low
+ 8.381010000e-07 V_low
+ 8.382000000e-07 V_low
+ 8.382010000e-07 V_low
+ 8.383000000e-07 V_low
+ 8.383010000e-07 V_low
+ 8.384000000e-07 V_low
+ 8.384010000e-07 V_low
+ 8.385000000e-07 V_low
+ 8.385010000e-07 V_low
+ 8.386000000e-07 V_low
+ 8.386010000e-07 V_low
+ 8.387000000e-07 V_low
+ 8.387010000e-07 V_low
+ 8.388000000e-07 V_low
+ 8.388010000e-07 V_low
+ 8.389000000e-07 V_low
+ 8.389010000e-07 V_low
+ 8.390000000e-07 V_low
+ 8.390010000e-07 V_low
+ 8.391000000e-07 V_low
+ 8.391010000e-07 V_low
+ 8.392000000e-07 V_low
+ 8.392010000e-07 V_low
+ 8.393000000e-07 V_low
+ 8.393010000e-07 V_low
+ 8.394000000e-07 V_low
+ 8.394010000e-07 V_low
+ 8.395000000e-07 V_low
+ 8.395010000e-07 V_low
+ 8.396000000e-07 V_low
+ 8.396010000e-07 V_low
+ 8.397000000e-07 V_low
+ 8.397010000e-07 V_low
+ 8.398000000e-07 V_low
+ 8.398010000e-07 V_low
+ 8.399000000e-07 V_low
+ 8.399010000e-07 V_low
+ 8.400000000e-07 V_low
+ 8.400010000e-07 V_low
+ 8.401000000e-07 V_low
+ 8.401010000e-07 V_low
+ 8.402000000e-07 V_low
+ 8.402010000e-07 V_low
+ 8.403000000e-07 V_low
+ 8.403010000e-07 V_low
+ 8.404000000e-07 V_low
+ 8.404010000e-07 V_low
+ 8.405000000e-07 V_low
+ 8.405010000e-07 V_low
+ 8.406000000e-07 V_low
+ 8.406010000e-07 V_low
+ 8.407000000e-07 V_low
+ 8.407010000e-07 V_low
+ 8.408000000e-07 V_low
+ 8.408010000e-07 V_low
+ 8.409000000e-07 V_low
+ 8.409010000e-07 V_low
+ 8.410000000e-07 V_low
+ 8.410010000e-07 V_low
+ 8.411000000e-07 V_low
+ 8.411010000e-07 V_low
+ 8.412000000e-07 V_low
+ 8.412010000e-07 V_low
+ 8.413000000e-07 V_low
+ 8.413010000e-07 V_low
+ 8.414000000e-07 V_low
+ 8.414010000e-07 V_low
+ 8.415000000e-07 V_low
+ 8.415010000e-07 V_low
+ 8.416000000e-07 V_low
+ 8.416010000e-07 V_low
+ 8.417000000e-07 V_low
+ 8.417010000e-07 V_low
+ 8.418000000e-07 V_low
+ 8.418010000e-07 V_low
+ 8.419000000e-07 V_low
+ 8.419010000e-07 V_hig
+ 8.420000000e-07 V_hig
+ 8.420010000e-07 V_hig
+ 8.421000000e-07 V_hig
+ 8.421010000e-07 V_hig
+ 8.422000000e-07 V_hig
+ 8.422010000e-07 V_hig
+ 8.423000000e-07 V_hig
+ 8.423010000e-07 V_hig
+ 8.424000000e-07 V_hig
+ 8.424010000e-07 V_hig
+ 8.425000000e-07 V_hig
+ 8.425010000e-07 V_hig
+ 8.426000000e-07 V_hig
+ 8.426010000e-07 V_hig
+ 8.427000000e-07 V_hig
+ 8.427010000e-07 V_hig
+ 8.428000000e-07 V_hig
+ 8.428010000e-07 V_hig
+ 8.429000000e-07 V_hig
+ 8.429010000e-07 V_hig
+ 8.430000000e-07 V_hig
+ 8.430010000e-07 V_hig
+ 8.431000000e-07 V_hig
+ 8.431010000e-07 V_hig
+ 8.432000000e-07 V_hig
+ 8.432010000e-07 V_hig
+ 8.433000000e-07 V_hig
+ 8.433010000e-07 V_hig
+ 8.434000000e-07 V_hig
+ 8.434010000e-07 V_hig
+ 8.435000000e-07 V_hig
+ 8.435010000e-07 V_hig
+ 8.436000000e-07 V_hig
+ 8.436010000e-07 V_hig
+ 8.437000000e-07 V_hig
+ 8.437010000e-07 V_hig
+ 8.438000000e-07 V_hig
+ 8.438010000e-07 V_hig
+ 8.439000000e-07 V_hig
+ 8.439010000e-07 V_hig
+ 8.440000000e-07 V_hig
+ 8.440010000e-07 V_hig
+ 8.441000000e-07 V_hig
+ 8.441010000e-07 V_hig
+ 8.442000000e-07 V_hig
+ 8.442010000e-07 V_hig
+ 8.443000000e-07 V_hig
+ 8.443010000e-07 V_hig
+ 8.444000000e-07 V_hig
+ 8.444010000e-07 V_hig
+ 8.445000000e-07 V_hig
+ 8.445010000e-07 V_hig
+ 8.446000000e-07 V_hig
+ 8.446010000e-07 V_hig
+ 8.447000000e-07 V_hig
+ 8.447010000e-07 V_hig
+ 8.448000000e-07 V_hig
+ 8.448010000e-07 V_hig
+ 8.449000000e-07 V_hig
+ 8.449010000e-07 V_hig
+ 8.450000000e-07 V_hig
+ 8.450010000e-07 V_hig
+ 8.451000000e-07 V_hig
+ 8.451010000e-07 V_hig
+ 8.452000000e-07 V_hig
+ 8.452010000e-07 V_hig
+ 8.453000000e-07 V_hig
+ 8.453010000e-07 V_hig
+ 8.454000000e-07 V_hig
+ 8.454010000e-07 V_hig
+ 8.455000000e-07 V_hig
+ 8.455010000e-07 V_hig
+ 8.456000000e-07 V_hig
+ 8.456010000e-07 V_hig
+ 8.457000000e-07 V_hig
+ 8.457010000e-07 V_hig
+ 8.458000000e-07 V_hig
+ 8.458010000e-07 V_hig
+ 8.459000000e-07 V_hig
+ 8.459010000e-07 V_hig
+ 8.460000000e-07 V_hig
+ 8.460010000e-07 V_hig
+ 8.461000000e-07 V_hig
+ 8.461010000e-07 V_hig
+ 8.462000000e-07 V_hig
+ 8.462010000e-07 V_hig
+ 8.463000000e-07 V_hig
+ 8.463010000e-07 V_hig
+ 8.464000000e-07 V_hig
+ 8.464010000e-07 V_hig
+ 8.465000000e-07 V_hig
+ 8.465010000e-07 V_hig
+ 8.466000000e-07 V_hig
+ 8.466010000e-07 V_hig
+ 8.467000000e-07 V_hig
+ 8.467010000e-07 V_hig
+ 8.468000000e-07 V_hig
+ 8.468010000e-07 V_hig
+ 8.469000000e-07 V_hig
+ 8.469010000e-07 V_hig
+ 8.470000000e-07 V_hig
+ 8.470010000e-07 V_hig
+ 8.471000000e-07 V_hig
+ 8.471010000e-07 V_hig
+ 8.472000000e-07 V_hig
+ 8.472010000e-07 V_hig
+ 8.473000000e-07 V_hig
+ 8.473010000e-07 V_hig
+ 8.474000000e-07 V_hig
+ 8.474010000e-07 V_hig
+ 8.475000000e-07 V_hig
+ 8.475010000e-07 V_hig
+ 8.476000000e-07 V_hig
+ 8.476010000e-07 V_hig
+ 8.477000000e-07 V_hig
+ 8.477010000e-07 V_hig
+ 8.478000000e-07 V_hig
+ 8.478010000e-07 V_hig
+ 8.479000000e-07 V_hig
+ 8.479010000e-07 V_hig
+ 8.480000000e-07 V_hig
+ 8.480010000e-07 V_hig
+ 8.481000000e-07 V_hig
+ 8.481010000e-07 V_hig
+ 8.482000000e-07 V_hig
+ 8.482010000e-07 V_hig
+ 8.483000000e-07 V_hig
+ 8.483010000e-07 V_hig
+ 8.484000000e-07 V_hig
+ 8.484010000e-07 V_hig
+ 8.485000000e-07 V_hig
+ 8.485010000e-07 V_hig
+ 8.486000000e-07 V_hig
+ 8.486010000e-07 V_hig
+ 8.487000000e-07 V_hig
+ 8.487010000e-07 V_hig
+ 8.488000000e-07 V_hig
+ 8.488010000e-07 V_hig
+ 8.489000000e-07 V_hig
+ 8.489010000e-07 V_low
+ 8.490000000e-07 V_low
+ 8.490010000e-07 V_low
+ 8.491000000e-07 V_low
+ 8.491010000e-07 V_low
+ 8.492000000e-07 V_low
+ 8.492010000e-07 V_low
+ 8.493000000e-07 V_low
+ 8.493010000e-07 V_low
+ 8.494000000e-07 V_low
+ 8.494010000e-07 V_low
+ 8.495000000e-07 V_low
+ 8.495010000e-07 V_low
+ 8.496000000e-07 V_low
+ 8.496010000e-07 V_low
+ 8.497000000e-07 V_low
+ 8.497010000e-07 V_low
+ 8.498000000e-07 V_low
+ 8.498010000e-07 V_low
+ 8.499000000e-07 V_low
+ 8.499010000e-07 V_hig
+ 8.500000000e-07 V_hig
+ 8.500010000e-07 V_hig
+ 8.501000000e-07 V_hig
+ 8.501010000e-07 V_hig
+ 8.502000000e-07 V_hig
+ 8.502010000e-07 V_hig
+ 8.503000000e-07 V_hig
+ 8.503010000e-07 V_hig
+ 8.504000000e-07 V_hig
+ 8.504010000e-07 V_hig
+ 8.505000000e-07 V_hig
+ 8.505010000e-07 V_hig
+ 8.506000000e-07 V_hig
+ 8.506010000e-07 V_hig
+ 8.507000000e-07 V_hig
+ 8.507010000e-07 V_hig
+ 8.508000000e-07 V_hig
+ 8.508010000e-07 V_hig
+ 8.509000000e-07 V_hig
+ 8.509010000e-07 V_hig
+ 8.510000000e-07 V_hig
+ 8.510010000e-07 V_hig
+ 8.511000000e-07 V_hig
+ 8.511010000e-07 V_hig
+ 8.512000000e-07 V_hig
+ 8.512010000e-07 V_hig
+ 8.513000000e-07 V_hig
+ 8.513010000e-07 V_hig
+ 8.514000000e-07 V_hig
+ 8.514010000e-07 V_hig
+ 8.515000000e-07 V_hig
+ 8.515010000e-07 V_hig
+ 8.516000000e-07 V_hig
+ 8.516010000e-07 V_hig
+ 8.517000000e-07 V_hig
+ 8.517010000e-07 V_hig
+ 8.518000000e-07 V_hig
+ 8.518010000e-07 V_hig
+ 8.519000000e-07 V_hig
+ 8.519010000e-07 V_hig
+ 8.520000000e-07 V_hig
+ 8.520010000e-07 V_hig
+ 8.521000000e-07 V_hig
+ 8.521010000e-07 V_hig
+ 8.522000000e-07 V_hig
+ 8.522010000e-07 V_hig
+ 8.523000000e-07 V_hig
+ 8.523010000e-07 V_hig
+ 8.524000000e-07 V_hig
+ 8.524010000e-07 V_hig
+ 8.525000000e-07 V_hig
+ 8.525010000e-07 V_hig
+ 8.526000000e-07 V_hig
+ 8.526010000e-07 V_hig
+ 8.527000000e-07 V_hig
+ 8.527010000e-07 V_hig
+ 8.528000000e-07 V_hig
+ 8.528010000e-07 V_hig
+ 8.529000000e-07 V_hig
+ 8.529010000e-07 V_low
+ 8.530000000e-07 V_low
+ 8.530010000e-07 V_low
+ 8.531000000e-07 V_low
+ 8.531010000e-07 V_low
+ 8.532000000e-07 V_low
+ 8.532010000e-07 V_low
+ 8.533000000e-07 V_low
+ 8.533010000e-07 V_low
+ 8.534000000e-07 V_low
+ 8.534010000e-07 V_low
+ 8.535000000e-07 V_low
+ 8.535010000e-07 V_low
+ 8.536000000e-07 V_low
+ 8.536010000e-07 V_low
+ 8.537000000e-07 V_low
+ 8.537010000e-07 V_low
+ 8.538000000e-07 V_low
+ 8.538010000e-07 V_low
+ 8.539000000e-07 V_low
+ 8.539010000e-07 V_low
+ 8.540000000e-07 V_low
+ 8.540010000e-07 V_low
+ 8.541000000e-07 V_low
+ 8.541010000e-07 V_low
+ 8.542000000e-07 V_low
+ 8.542010000e-07 V_low
+ 8.543000000e-07 V_low
+ 8.543010000e-07 V_low
+ 8.544000000e-07 V_low
+ 8.544010000e-07 V_low
+ 8.545000000e-07 V_low
+ 8.545010000e-07 V_low
+ 8.546000000e-07 V_low
+ 8.546010000e-07 V_low
+ 8.547000000e-07 V_low
+ 8.547010000e-07 V_low
+ 8.548000000e-07 V_low
+ 8.548010000e-07 V_low
+ 8.549000000e-07 V_low
+ 8.549010000e-07 V_low
+ 8.550000000e-07 V_low
+ 8.550010000e-07 V_low
+ 8.551000000e-07 V_low
+ 8.551010000e-07 V_low
+ 8.552000000e-07 V_low
+ 8.552010000e-07 V_low
+ 8.553000000e-07 V_low
+ 8.553010000e-07 V_low
+ 8.554000000e-07 V_low
+ 8.554010000e-07 V_low
+ 8.555000000e-07 V_low
+ 8.555010000e-07 V_low
+ 8.556000000e-07 V_low
+ 8.556010000e-07 V_low
+ 8.557000000e-07 V_low
+ 8.557010000e-07 V_low
+ 8.558000000e-07 V_low
+ 8.558010000e-07 V_low
+ 8.559000000e-07 V_low
+ 8.559010000e-07 V_low
+ 8.560000000e-07 V_low
+ 8.560010000e-07 V_low
+ 8.561000000e-07 V_low
+ 8.561010000e-07 V_low
+ 8.562000000e-07 V_low
+ 8.562010000e-07 V_low
+ 8.563000000e-07 V_low
+ 8.563010000e-07 V_low
+ 8.564000000e-07 V_low
+ 8.564010000e-07 V_low
+ 8.565000000e-07 V_low
+ 8.565010000e-07 V_low
+ 8.566000000e-07 V_low
+ 8.566010000e-07 V_low
+ 8.567000000e-07 V_low
+ 8.567010000e-07 V_low
+ 8.568000000e-07 V_low
+ 8.568010000e-07 V_low
+ 8.569000000e-07 V_low
+ 8.569010000e-07 V_hig
+ 8.570000000e-07 V_hig
+ 8.570010000e-07 V_hig
+ 8.571000000e-07 V_hig
+ 8.571010000e-07 V_hig
+ 8.572000000e-07 V_hig
+ 8.572010000e-07 V_hig
+ 8.573000000e-07 V_hig
+ 8.573010000e-07 V_hig
+ 8.574000000e-07 V_hig
+ 8.574010000e-07 V_hig
+ 8.575000000e-07 V_hig
+ 8.575010000e-07 V_hig
+ 8.576000000e-07 V_hig
+ 8.576010000e-07 V_hig
+ 8.577000000e-07 V_hig
+ 8.577010000e-07 V_hig
+ 8.578000000e-07 V_hig
+ 8.578010000e-07 V_hig
+ 8.579000000e-07 V_hig
+ 8.579010000e-07 V_low
+ 8.580000000e-07 V_low
+ 8.580010000e-07 V_low
+ 8.581000000e-07 V_low
+ 8.581010000e-07 V_low
+ 8.582000000e-07 V_low
+ 8.582010000e-07 V_low
+ 8.583000000e-07 V_low
+ 8.583010000e-07 V_low
+ 8.584000000e-07 V_low
+ 8.584010000e-07 V_low
+ 8.585000000e-07 V_low
+ 8.585010000e-07 V_low
+ 8.586000000e-07 V_low
+ 8.586010000e-07 V_low
+ 8.587000000e-07 V_low
+ 8.587010000e-07 V_low
+ 8.588000000e-07 V_low
+ 8.588010000e-07 V_low
+ 8.589000000e-07 V_low
+ 8.589010000e-07 V_hig
+ 8.590000000e-07 V_hig
+ 8.590010000e-07 V_hig
+ 8.591000000e-07 V_hig
+ 8.591010000e-07 V_hig
+ 8.592000000e-07 V_hig
+ 8.592010000e-07 V_hig
+ 8.593000000e-07 V_hig
+ 8.593010000e-07 V_hig
+ 8.594000000e-07 V_hig
+ 8.594010000e-07 V_hig
+ 8.595000000e-07 V_hig
+ 8.595010000e-07 V_hig
+ 8.596000000e-07 V_hig
+ 8.596010000e-07 V_hig
+ 8.597000000e-07 V_hig
+ 8.597010000e-07 V_hig
+ 8.598000000e-07 V_hig
+ 8.598010000e-07 V_hig
+ 8.599000000e-07 V_hig
+ 8.599010000e-07 V_low
+ 8.600000000e-07 V_low
+ 8.600010000e-07 V_low
+ 8.601000000e-07 V_low
+ 8.601010000e-07 V_low
+ 8.602000000e-07 V_low
+ 8.602010000e-07 V_low
+ 8.603000000e-07 V_low
+ 8.603010000e-07 V_low
+ 8.604000000e-07 V_low
+ 8.604010000e-07 V_low
+ 8.605000000e-07 V_low
+ 8.605010000e-07 V_low
+ 8.606000000e-07 V_low
+ 8.606010000e-07 V_low
+ 8.607000000e-07 V_low
+ 8.607010000e-07 V_low
+ 8.608000000e-07 V_low
+ 8.608010000e-07 V_low
+ 8.609000000e-07 V_low
+ 8.609010000e-07 V_low
+ 8.610000000e-07 V_low
+ 8.610010000e-07 V_low
+ 8.611000000e-07 V_low
+ 8.611010000e-07 V_low
+ 8.612000000e-07 V_low
+ 8.612010000e-07 V_low
+ 8.613000000e-07 V_low
+ 8.613010000e-07 V_low
+ 8.614000000e-07 V_low
+ 8.614010000e-07 V_low
+ 8.615000000e-07 V_low
+ 8.615010000e-07 V_low
+ 8.616000000e-07 V_low
+ 8.616010000e-07 V_low
+ 8.617000000e-07 V_low
+ 8.617010000e-07 V_low
+ 8.618000000e-07 V_low
+ 8.618010000e-07 V_low
+ 8.619000000e-07 V_low
+ 8.619010000e-07 V_hig
+ 8.620000000e-07 V_hig
+ 8.620010000e-07 V_hig
+ 8.621000000e-07 V_hig
+ 8.621010000e-07 V_hig
+ 8.622000000e-07 V_hig
+ 8.622010000e-07 V_hig
+ 8.623000000e-07 V_hig
+ 8.623010000e-07 V_hig
+ 8.624000000e-07 V_hig
+ 8.624010000e-07 V_hig
+ 8.625000000e-07 V_hig
+ 8.625010000e-07 V_hig
+ 8.626000000e-07 V_hig
+ 8.626010000e-07 V_hig
+ 8.627000000e-07 V_hig
+ 8.627010000e-07 V_hig
+ 8.628000000e-07 V_hig
+ 8.628010000e-07 V_hig
+ 8.629000000e-07 V_hig
+ 8.629010000e-07 V_hig
+ 8.630000000e-07 V_hig
+ 8.630010000e-07 V_hig
+ 8.631000000e-07 V_hig
+ 8.631010000e-07 V_hig
+ 8.632000000e-07 V_hig
+ 8.632010000e-07 V_hig
+ 8.633000000e-07 V_hig
+ 8.633010000e-07 V_hig
+ 8.634000000e-07 V_hig
+ 8.634010000e-07 V_hig
+ 8.635000000e-07 V_hig
+ 8.635010000e-07 V_hig
+ 8.636000000e-07 V_hig
+ 8.636010000e-07 V_hig
+ 8.637000000e-07 V_hig
+ 8.637010000e-07 V_hig
+ 8.638000000e-07 V_hig
+ 8.638010000e-07 V_hig
+ 8.639000000e-07 V_hig
+ 8.639010000e-07 V_hig
+ 8.640000000e-07 V_hig
+ 8.640010000e-07 V_hig
+ 8.641000000e-07 V_hig
+ 8.641010000e-07 V_hig
+ 8.642000000e-07 V_hig
+ 8.642010000e-07 V_hig
+ 8.643000000e-07 V_hig
+ 8.643010000e-07 V_hig
+ 8.644000000e-07 V_hig
+ 8.644010000e-07 V_hig
+ 8.645000000e-07 V_hig
+ 8.645010000e-07 V_hig
+ 8.646000000e-07 V_hig
+ 8.646010000e-07 V_hig
+ 8.647000000e-07 V_hig
+ 8.647010000e-07 V_hig
+ 8.648000000e-07 V_hig
+ 8.648010000e-07 V_hig
+ 8.649000000e-07 V_hig
+ 8.649010000e-07 V_low
+ 8.650000000e-07 V_low
+ 8.650010000e-07 V_low
+ 8.651000000e-07 V_low
+ 8.651010000e-07 V_low
+ 8.652000000e-07 V_low
+ 8.652010000e-07 V_low
+ 8.653000000e-07 V_low
+ 8.653010000e-07 V_low
+ 8.654000000e-07 V_low
+ 8.654010000e-07 V_low
+ 8.655000000e-07 V_low
+ 8.655010000e-07 V_low
+ 8.656000000e-07 V_low
+ 8.656010000e-07 V_low
+ 8.657000000e-07 V_low
+ 8.657010000e-07 V_low
+ 8.658000000e-07 V_low
+ 8.658010000e-07 V_low
+ 8.659000000e-07 V_low
+ 8.659010000e-07 V_low
+ 8.660000000e-07 V_low
+ 8.660010000e-07 V_low
+ 8.661000000e-07 V_low
+ 8.661010000e-07 V_low
+ 8.662000000e-07 V_low
+ 8.662010000e-07 V_low
+ 8.663000000e-07 V_low
+ 8.663010000e-07 V_low
+ 8.664000000e-07 V_low
+ 8.664010000e-07 V_low
+ 8.665000000e-07 V_low
+ 8.665010000e-07 V_low
+ 8.666000000e-07 V_low
+ 8.666010000e-07 V_low
+ 8.667000000e-07 V_low
+ 8.667010000e-07 V_low
+ 8.668000000e-07 V_low
+ 8.668010000e-07 V_low
+ 8.669000000e-07 V_low
+ 8.669010000e-07 V_hig
+ 8.670000000e-07 V_hig
+ 8.670010000e-07 V_hig
+ 8.671000000e-07 V_hig
+ 8.671010000e-07 V_hig
+ 8.672000000e-07 V_hig
+ 8.672010000e-07 V_hig
+ 8.673000000e-07 V_hig
+ 8.673010000e-07 V_hig
+ 8.674000000e-07 V_hig
+ 8.674010000e-07 V_hig
+ 8.675000000e-07 V_hig
+ 8.675010000e-07 V_hig
+ 8.676000000e-07 V_hig
+ 8.676010000e-07 V_hig
+ 8.677000000e-07 V_hig
+ 8.677010000e-07 V_hig
+ 8.678000000e-07 V_hig
+ 8.678010000e-07 V_hig
+ 8.679000000e-07 V_hig
+ 8.679010000e-07 V_hig
+ 8.680000000e-07 V_hig
+ 8.680010000e-07 V_hig
+ 8.681000000e-07 V_hig
+ 8.681010000e-07 V_hig
+ 8.682000000e-07 V_hig
+ 8.682010000e-07 V_hig
+ 8.683000000e-07 V_hig
+ 8.683010000e-07 V_hig
+ 8.684000000e-07 V_hig
+ 8.684010000e-07 V_hig
+ 8.685000000e-07 V_hig
+ 8.685010000e-07 V_hig
+ 8.686000000e-07 V_hig
+ 8.686010000e-07 V_hig
+ 8.687000000e-07 V_hig
+ 8.687010000e-07 V_hig
+ 8.688000000e-07 V_hig
+ 8.688010000e-07 V_hig
+ 8.689000000e-07 V_hig
+ 8.689010000e-07 V_hig
+ 8.690000000e-07 V_hig
+ 8.690010000e-07 V_hig
+ 8.691000000e-07 V_hig
+ 8.691010000e-07 V_hig
+ 8.692000000e-07 V_hig
+ 8.692010000e-07 V_hig
+ 8.693000000e-07 V_hig
+ 8.693010000e-07 V_hig
+ 8.694000000e-07 V_hig
+ 8.694010000e-07 V_hig
+ 8.695000000e-07 V_hig
+ 8.695010000e-07 V_hig
+ 8.696000000e-07 V_hig
+ 8.696010000e-07 V_hig
+ 8.697000000e-07 V_hig
+ 8.697010000e-07 V_hig
+ 8.698000000e-07 V_hig
+ 8.698010000e-07 V_hig
+ 8.699000000e-07 V_hig
+ 8.699010000e-07 V_low
+ 8.700000000e-07 V_low
+ 8.700010000e-07 V_low
+ 8.701000000e-07 V_low
+ 8.701010000e-07 V_low
+ 8.702000000e-07 V_low
+ 8.702010000e-07 V_low
+ 8.703000000e-07 V_low
+ 8.703010000e-07 V_low
+ 8.704000000e-07 V_low
+ 8.704010000e-07 V_low
+ 8.705000000e-07 V_low
+ 8.705010000e-07 V_low
+ 8.706000000e-07 V_low
+ 8.706010000e-07 V_low
+ 8.707000000e-07 V_low
+ 8.707010000e-07 V_low
+ 8.708000000e-07 V_low
+ 8.708010000e-07 V_low
+ 8.709000000e-07 V_low
+ 8.709010000e-07 V_low
+ 8.710000000e-07 V_low
+ 8.710010000e-07 V_low
+ 8.711000000e-07 V_low
+ 8.711010000e-07 V_low
+ 8.712000000e-07 V_low
+ 8.712010000e-07 V_low
+ 8.713000000e-07 V_low
+ 8.713010000e-07 V_low
+ 8.714000000e-07 V_low
+ 8.714010000e-07 V_low
+ 8.715000000e-07 V_low
+ 8.715010000e-07 V_low
+ 8.716000000e-07 V_low
+ 8.716010000e-07 V_low
+ 8.717000000e-07 V_low
+ 8.717010000e-07 V_low
+ 8.718000000e-07 V_low
+ 8.718010000e-07 V_low
+ 8.719000000e-07 V_low
+ 8.719010000e-07 V_hig
+ 8.720000000e-07 V_hig
+ 8.720010000e-07 V_hig
+ 8.721000000e-07 V_hig
+ 8.721010000e-07 V_hig
+ 8.722000000e-07 V_hig
+ 8.722010000e-07 V_hig
+ 8.723000000e-07 V_hig
+ 8.723010000e-07 V_hig
+ 8.724000000e-07 V_hig
+ 8.724010000e-07 V_hig
+ 8.725000000e-07 V_hig
+ 8.725010000e-07 V_hig
+ 8.726000000e-07 V_hig
+ 8.726010000e-07 V_hig
+ 8.727000000e-07 V_hig
+ 8.727010000e-07 V_hig
+ 8.728000000e-07 V_hig
+ 8.728010000e-07 V_hig
+ 8.729000000e-07 V_hig
+ 8.729010000e-07 V_low
+ 8.730000000e-07 V_low
+ 8.730010000e-07 V_low
+ 8.731000000e-07 V_low
+ 8.731010000e-07 V_low
+ 8.732000000e-07 V_low
+ 8.732010000e-07 V_low
+ 8.733000000e-07 V_low
+ 8.733010000e-07 V_low
+ 8.734000000e-07 V_low
+ 8.734010000e-07 V_low
+ 8.735000000e-07 V_low
+ 8.735010000e-07 V_low
+ 8.736000000e-07 V_low
+ 8.736010000e-07 V_low
+ 8.737000000e-07 V_low
+ 8.737010000e-07 V_low
+ 8.738000000e-07 V_low
+ 8.738010000e-07 V_low
+ 8.739000000e-07 V_low
+ 8.739010000e-07 V_low
+ 8.740000000e-07 V_low
+ 8.740010000e-07 V_low
+ 8.741000000e-07 V_low
+ 8.741010000e-07 V_low
+ 8.742000000e-07 V_low
+ 8.742010000e-07 V_low
+ 8.743000000e-07 V_low
+ 8.743010000e-07 V_low
+ 8.744000000e-07 V_low
+ 8.744010000e-07 V_low
+ 8.745000000e-07 V_low
+ 8.745010000e-07 V_low
+ 8.746000000e-07 V_low
+ 8.746010000e-07 V_low
+ 8.747000000e-07 V_low
+ 8.747010000e-07 V_low
+ 8.748000000e-07 V_low
+ 8.748010000e-07 V_low
+ 8.749000000e-07 V_low
+ 8.749010000e-07 V_low
+ 8.750000000e-07 V_low
+ 8.750010000e-07 V_low
+ 8.751000000e-07 V_low
+ 8.751010000e-07 V_low
+ 8.752000000e-07 V_low
+ 8.752010000e-07 V_low
+ 8.753000000e-07 V_low
+ 8.753010000e-07 V_low
+ 8.754000000e-07 V_low
+ 8.754010000e-07 V_low
+ 8.755000000e-07 V_low
+ 8.755010000e-07 V_low
+ 8.756000000e-07 V_low
+ 8.756010000e-07 V_low
+ 8.757000000e-07 V_low
+ 8.757010000e-07 V_low
+ 8.758000000e-07 V_low
+ 8.758010000e-07 V_low
+ 8.759000000e-07 V_low
+ 8.759010000e-07 V_hig
+ 8.760000000e-07 V_hig
+ 8.760010000e-07 V_hig
+ 8.761000000e-07 V_hig
+ 8.761010000e-07 V_hig
+ 8.762000000e-07 V_hig
+ 8.762010000e-07 V_hig
+ 8.763000000e-07 V_hig
+ 8.763010000e-07 V_hig
+ 8.764000000e-07 V_hig
+ 8.764010000e-07 V_hig
+ 8.765000000e-07 V_hig
+ 8.765010000e-07 V_hig
+ 8.766000000e-07 V_hig
+ 8.766010000e-07 V_hig
+ 8.767000000e-07 V_hig
+ 8.767010000e-07 V_hig
+ 8.768000000e-07 V_hig
+ 8.768010000e-07 V_hig
+ 8.769000000e-07 V_hig
+ 8.769010000e-07 V_hig
+ 8.770000000e-07 V_hig
+ 8.770010000e-07 V_hig
+ 8.771000000e-07 V_hig
+ 8.771010000e-07 V_hig
+ 8.772000000e-07 V_hig
+ 8.772010000e-07 V_hig
+ 8.773000000e-07 V_hig
+ 8.773010000e-07 V_hig
+ 8.774000000e-07 V_hig
+ 8.774010000e-07 V_hig
+ 8.775000000e-07 V_hig
+ 8.775010000e-07 V_hig
+ 8.776000000e-07 V_hig
+ 8.776010000e-07 V_hig
+ 8.777000000e-07 V_hig
+ 8.777010000e-07 V_hig
+ 8.778000000e-07 V_hig
+ 8.778010000e-07 V_hig
+ 8.779000000e-07 V_hig
+ 8.779010000e-07 V_low
+ 8.780000000e-07 V_low
+ 8.780010000e-07 V_low
+ 8.781000000e-07 V_low
+ 8.781010000e-07 V_low
+ 8.782000000e-07 V_low
+ 8.782010000e-07 V_low
+ 8.783000000e-07 V_low
+ 8.783010000e-07 V_low
+ 8.784000000e-07 V_low
+ 8.784010000e-07 V_low
+ 8.785000000e-07 V_low
+ 8.785010000e-07 V_low
+ 8.786000000e-07 V_low
+ 8.786010000e-07 V_low
+ 8.787000000e-07 V_low
+ 8.787010000e-07 V_low
+ 8.788000000e-07 V_low
+ 8.788010000e-07 V_low
+ 8.789000000e-07 V_low
+ 8.789010000e-07 V_low
+ 8.790000000e-07 V_low
+ 8.790010000e-07 V_low
+ 8.791000000e-07 V_low
+ 8.791010000e-07 V_low
+ 8.792000000e-07 V_low
+ 8.792010000e-07 V_low
+ 8.793000000e-07 V_low
+ 8.793010000e-07 V_low
+ 8.794000000e-07 V_low
+ 8.794010000e-07 V_low
+ 8.795000000e-07 V_low
+ 8.795010000e-07 V_low
+ 8.796000000e-07 V_low
+ 8.796010000e-07 V_low
+ 8.797000000e-07 V_low
+ 8.797010000e-07 V_low
+ 8.798000000e-07 V_low
+ 8.798010000e-07 V_low
+ 8.799000000e-07 V_low
+ 8.799010000e-07 V_hig
+ 8.800000000e-07 V_hig
+ 8.800010000e-07 V_hig
+ 8.801000000e-07 V_hig
+ 8.801010000e-07 V_hig
+ 8.802000000e-07 V_hig
+ 8.802010000e-07 V_hig
+ 8.803000000e-07 V_hig
+ 8.803010000e-07 V_hig
+ 8.804000000e-07 V_hig
+ 8.804010000e-07 V_hig
+ 8.805000000e-07 V_hig
+ 8.805010000e-07 V_hig
+ 8.806000000e-07 V_hig
+ 8.806010000e-07 V_hig
+ 8.807000000e-07 V_hig
+ 8.807010000e-07 V_hig
+ 8.808000000e-07 V_hig
+ 8.808010000e-07 V_hig
+ 8.809000000e-07 V_hig
+ 8.809010000e-07 V_low
+ 8.810000000e-07 V_low
+ 8.810010000e-07 V_low
+ 8.811000000e-07 V_low
+ 8.811010000e-07 V_low
+ 8.812000000e-07 V_low
+ 8.812010000e-07 V_low
+ 8.813000000e-07 V_low
+ 8.813010000e-07 V_low
+ 8.814000000e-07 V_low
+ 8.814010000e-07 V_low
+ 8.815000000e-07 V_low
+ 8.815010000e-07 V_low
+ 8.816000000e-07 V_low
+ 8.816010000e-07 V_low
+ 8.817000000e-07 V_low
+ 8.817010000e-07 V_low
+ 8.818000000e-07 V_low
+ 8.818010000e-07 V_low
+ 8.819000000e-07 V_low
+ 8.819010000e-07 V_hig
+ 8.820000000e-07 V_hig
+ 8.820010000e-07 V_hig
+ 8.821000000e-07 V_hig
+ 8.821010000e-07 V_hig
+ 8.822000000e-07 V_hig
+ 8.822010000e-07 V_hig
+ 8.823000000e-07 V_hig
+ 8.823010000e-07 V_hig
+ 8.824000000e-07 V_hig
+ 8.824010000e-07 V_hig
+ 8.825000000e-07 V_hig
+ 8.825010000e-07 V_hig
+ 8.826000000e-07 V_hig
+ 8.826010000e-07 V_hig
+ 8.827000000e-07 V_hig
+ 8.827010000e-07 V_hig
+ 8.828000000e-07 V_hig
+ 8.828010000e-07 V_hig
+ 8.829000000e-07 V_hig
+ 8.829010000e-07 V_hig
+ 8.830000000e-07 V_hig
+ 8.830010000e-07 V_hig
+ 8.831000000e-07 V_hig
+ 8.831010000e-07 V_hig
+ 8.832000000e-07 V_hig
+ 8.832010000e-07 V_hig
+ 8.833000000e-07 V_hig
+ 8.833010000e-07 V_hig
+ 8.834000000e-07 V_hig
+ 8.834010000e-07 V_hig
+ 8.835000000e-07 V_hig
+ 8.835010000e-07 V_hig
+ 8.836000000e-07 V_hig
+ 8.836010000e-07 V_hig
+ 8.837000000e-07 V_hig
+ 8.837010000e-07 V_hig
+ 8.838000000e-07 V_hig
+ 8.838010000e-07 V_hig
+ 8.839000000e-07 V_hig
+ 8.839010000e-07 V_low
+ 8.840000000e-07 V_low
+ 8.840010000e-07 V_low
+ 8.841000000e-07 V_low
+ 8.841010000e-07 V_low
+ 8.842000000e-07 V_low
+ 8.842010000e-07 V_low
+ 8.843000000e-07 V_low
+ 8.843010000e-07 V_low
+ 8.844000000e-07 V_low
+ 8.844010000e-07 V_low
+ 8.845000000e-07 V_low
+ 8.845010000e-07 V_low
+ 8.846000000e-07 V_low
+ 8.846010000e-07 V_low
+ 8.847000000e-07 V_low
+ 8.847010000e-07 V_low
+ 8.848000000e-07 V_low
+ 8.848010000e-07 V_low
+ 8.849000000e-07 V_low
+ 8.849010000e-07 V_low
+ 8.850000000e-07 V_low
+ 8.850010000e-07 V_low
+ 8.851000000e-07 V_low
+ 8.851010000e-07 V_low
+ 8.852000000e-07 V_low
+ 8.852010000e-07 V_low
+ 8.853000000e-07 V_low
+ 8.853010000e-07 V_low
+ 8.854000000e-07 V_low
+ 8.854010000e-07 V_low
+ 8.855000000e-07 V_low
+ 8.855010000e-07 V_low
+ 8.856000000e-07 V_low
+ 8.856010000e-07 V_low
+ 8.857000000e-07 V_low
+ 8.857010000e-07 V_low
+ 8.858000000e-07 V_low
+ 8.858010000e-07 V_low
+ 8.859000000e-07 V_low
+ 8.859010000e-07 V_low
+ 8.860000000e-07 V_low
+ 8.860010000e-07 V_low
+ 8.861000000e-07 V_low
+ 8.861010000e-07 V_low
+ 8.862000000e-07 V_low
+ 8.862010000e-07 V_low
+ 8.863000000e-07 V_low
+ 8.863010000e-07 V_low
+ 8.864000000e-07 V_low
+ 8.864010000e-07 V_low
+ 8.865000000e-07 V_low
+ 8.865010000e-07 V_low
+ 8.866000000e-07 V_low
+ 8.866010000e-07 V_low
+ 8.867000000e-07 V_low
+ 8.867010000e-07 V_low
+ 8.868000000e-07 V_low
+ 8.868010000e-07 V_low
+ 8.869000000e-07 V_low
+ 8.869010000e-07 V_low
+ 8.870000000e-07 V_low
+ 8.870010000e-07 V_low
+ 8.871000000e-07 V_low
+ 8.871010000e-07 V_low
+ 8.872000000e-07 V_low
+ 8.872010000e-07 V_low
+ 8.873000000e-07 V_low
+ 8.873010000e-07 V_low
+ 8.874000000e-07 V_low
+ 8.874010000e-07 V_low
+ 8.875000000e-07 V_low
+ 8.875010000e-07 V_low
+ 8.876000000e-07 V_low
+ 8.876010000e-07 V_low
+ 8.877000000e-07 V_low
+ 8.877010000e-07 V_low
+ 8.878000000e-07 V_low
+ 8.878010000e-07 V_low
+ 8.879000000e-07 V_low
+ 8.879010000e-07 V_low
+ 8.880000000e-07 V_low
+ 8.880010000e-07 V_low
+ 8.881000000e-07 V_low
+ 8.881010000e-07 V_low
+ 8.882000000e-07 V_low
+ 8.882010000e-07 V_low
+ 8.883000000e-07 V_low
+ 8.883010000e-07 V_low
+ 8.884000000e-07 V_low
+ 8.884010000e-07 V_low
+ 8.885000000e-07 V_low
+ 8.885010000e-07 V_low
+ 8.886000000e-07 V_low
+ 8.886010000e-07 V_low
+ 8.887000000e-07 V_low
+ 8.887010000e-07 V_low
+ 8.888000000e-07 V_low
+ 8.888010000e-07 V_low
+ 8.889000000e-07 V_low
+ 8.889010000e-07 V_hig
+ 8.890000000e-07 V_hig
+ 8.890010000e-07 V_hig
+ 8.891000000e-07 V_hig
+ 8.891010000e-07 V_hig
+ 8.892000000e-07 V_hig
+ 8.892010000e-07 V_hig
+ 8.893000000e-07 V_hig
+ 8.893010000e-07 V_hig
+ 8.894000000e-07 V_hig
+ 8.894010000e-07 V_hig
+ 8.895000000e-07 V_hig
+ 8.895010000e-07 V_hig
+ 8.896000000e-07 V_hig
+ 8.896010000e-07 V_hig
+ 8.897000000e-07 V_hig
+ 8.897010000e-07 V_hig
+ 8.898000000e-07 V_hig
+ 8.898010000e-07 V_hig
+ 8.899000000e-07 V_hig
+ 8.899010000e-07 V_hig
+ 8.900000000e-07 V_hig
+ 8.900010000e-07 V_hig
+ 8.901000000e-07 V_hig
+ 8.901010000e-07 V_hig
+ 8.902000000e-07 V_hig
+ 8.902010000e-07 V_hig
+ 8.903000000e-07 V_hig
+ 8.903010000e-07 V_hig
+ 8.904000000e-07 V_hig
+ 8.904010000e-07 V_hig
+ 8.905000000e-07 V_hig
+ 8.905010000e-07 V_hig
+ 8.906000000e-07 V_hig
+ 8.906010000e-07 V_hig
+ 8.907000000e-07 V_hig
+ 8.907010000e-07 V_hig
+ 8.908000000e-07 V_hig
+ 8.908010000e-07 V_hig
+ 8.909000000e-07 V_hig
+ 8.909010000e-07 V_hig
+ 8.910000000e-07 V_hig
+ 8.910010000e-07 V_hig
+ 8.911000000e-07 V_hig
+ 8.911010000e-07 V_hig
+ 8.912000000e-07 V_hig
+ 8.912010000e-07 V_hig
+ 8.913000000e-07 V_hig
+ 8.913010000e-07 V_hig
+ 8.914000000e-07 V_hig
+ 8.914010000e-07 V_hig
+ 8.915000000e-07 V_hig
+ 8.915010000e-07 V_hig
+ 8.916000000e-07 V_hig
+ 8.916010000e-07 V_hig
+ 8.917000000e-07 V_hig
+ 8.917010000e-07 V_hig
+ 8.918000000e-07 V_hig
+ 8.918010000e-07 V_hig
+ 8.919000000e-07 V_hig
+ 8.919010000e-07 V_low
+ 8.920000000e-07 V_low
+ 8.920010000e-07 V_low
+ 8.921000000e-07 V_low
+ 8.921010000e-07 V_low
+ 8.922000000e-07 V_low
+ 8.922010000e-07 V_low
+ 8.923000000e-07 V_low
+ 8.923010000e-07 V_low
+ 8.924000000e-07 V_low
+ 8.924010000e-07 V_low
+ 8.925000000e-07 V_low
+ 8.925010000e-07 V_low
+ 8.926000000e-07 V_low
+ 8.926010000e-07 V_low
+ 8.927000000e-07 V_low
+ 8.927010000e-07 V_low
+ 8.928000000e-07 V_low
+ 8.928010000e-07 V_low
+ 8.929000000e-07 V_low
+ 8.929010000e-07 V_hig
+ 8.930000000e-07 V_hig
+ 8.930010000e-07 V_hig
+ 8.931000000e-07 V_hig
+ 8.931010000e-07 V_hig
+ 8.932000000e-07 V_hig
+ 8.932010000e-07 V_hig
+ 8.933000000e-07 V_hig
+ 8.933010000e-07 V_hig
+ 8.934000000e-07 V_hig
+ 8.934010000e-07 V_hig
+ 8.935000000e-07 V_hig
+ 8.935010000e-07 V_hig
+ 8.936000000e-07 V_hig
+ 8.936010000e-07 V_hig
+ 8.937000000e-07 V_hig
+ 8.937010000e-07 V_hig
+ 8.938000000e-07 V_hig
+ 8.938010000e-07 V_hig
+ 8.939000000e-07 V_hig
+ 8.939010000e-07 V_low
+ 8.940000000e-07 V_low
+ 8.940010000e-07 V_low
+ 8.941000000e-07 V_low
+ 8.941010000e-07 V_low
+ 8.942000000e-07 V_low
+ 8.942010000e-07 V_low
+ 8.943000000e-07 V_low
+ 8.943010000e-07 V_low
+ 8.944000000e-07 V_low
+ 8.944010000e-07 V_low
+ 8.945000000e-07 V_low
+ 8.945010000e-07 V_low
+ 8.946000000e-07 V_low
+ 8.946010000e-07 V_low
+ 8.947000000e-07 V_low
+ 8.947010000e-07 V_low
+ 8.948000000e-07 V_low
+ 8.948010000e-07 V_low
+ 8.949000000e-07 V_low
+ 8.949010000e-07 V_hig
+ 8.950000000e-07 V_hig
+ 8.950010000e-07 V_hig
+ 8.951000000e-07 V_hig
+ 8.951010000e-07 V_hig
+ 8.952000000e-07 V_hig
+ 8.952010000e-07 V_hig
+ 8.953000000e-07 V_hig
+ 8.953010000e-07 V_hig
+ 8.954000000e-07 V_hig
+ 8.954010000e-07 V_hig
+ 8.955000000e-07 V_hig
+ 8.955010000e-07 V_hig
+ 8.956000000e-07 V_hig
+ 8.956010000e-07 V_hig
+ 8.957000000e-07 V_hig
+ 8.957010000e-07 V_hig
+ 8.958000000e-07 V_hig
+ 8.958010000e-07 V_hig
+ 8.959000000e-07 V_hig
+ 8.959010000e-07 V_low
+ 8.960000000e-07 V_low
+ 8.960010000e-07 V_low
+ 8.961000000e-07 V_low
+ 8.961010000e-07 V_low
+ 8.962000000e-07 V_low
+ 8.962010000e-07 V_low
+ 8.963000000e-07 V_low
+ 8.963010000e-07 V_low
+ 8.964000000e-07 V_low
+ 8.964010000e-07 V_low
+ 8.965000000e-07 V_low
+ 8.965010000e-07 V_low
+ 8.966000000e-07 V_low
+ 8.966010000e-07 V_low
+ 8.967000000e-07 V_low
+ 8.967010000e-07 V_low
+ 8.968000000e-07 V_low
+ 8.968010000e-07 V_low
+ 8.969000000e-07 V_low
+ 8.969010000e-07 V_low
+ 8.970000000e-07 V_low
+ 8.970010000e-07 V_low
+ 8.971000000e-07 V_low
+ 8.971010000e-07 V_low
+ 8.972000000e-07 V_low
+ 8.972010000e-07 V_low
+ 8.973000000e-07 V_low
+ 8.973010000e-07 V_low
+ 8.974000000e-07 V_low
+ 8.974010000e-07 V_low
+ 8.975000000e-07 V_low
+ 8.975010000e-07 V_low
+ 8.976000000e-07 V_low
+ 8.976010000e-07 V_low
+ 8.977000000e-07 V_low
+ 8.977010000e-07 V_low
+ 8.978000000e-07 V_low
+ 8.978010000e-07 V_low
+ 8.979000000e-07 V_low
+ 8.979010000e-07 V_hig
+ 8.980000000e-07 V_hig
+ 8.980010000e-07 V_hig
+ 8.981000000e-07 V_hig
+ 8.981010000e-07 V_hig
+ 8.982000000e-07 V_hig
+ 8.982010000e-07 V_hig
+ 8.983000000e-07 V_hig
+ 8.983010000e-07 V_hig
+ 8.984000000e-07 V_hig
+ 8.984010000e-07 V_hig
+ 8.985000000e-07 V_hig
+ 8.985010000e-07 V_hig
+ 8.986000000e-07 V_hig
+ 8.986010000e-07 V_hig
+ 8.987000000e-07 V_hig
+ 8.987010000e-07 V_hig
+ 8.988000000e-07 V_hig
+ 8.988010000e-07 V_hig
+ 8.989000000e-07 V_hig
+ 8.989010000e-07 V_hig
+ 8.990000000e-07 V_hig
+ 8.990010000e-07 V_hig
+ 8.991000000e-07 V_hig
+ 8.991010000e-07 V_hig
+ 8.992000000e-07 V_hig
+ 8.992010000e-07 V_hig
+ 8.993000000e-07 V_hig
+ 8.993010000e-07 V_hig
+ 8.994000000e-07 V_hig
+ 8.994010000e-07 V_hig
+ 8.995000000e-07 V_hig
+ 8.995010000e-07 V_hig
+ 8.996000000e-07 V_hig
+ 8.996010000e-07 V_hig
+ 8.997000000e-07 V_hig
+ 8.997010000e-07 V_hig
+ 8.998000000e-07 V_hig
+ 8.998010000e-07 V_hig
+ 8.999000000e-07 V_hig
+ 8.999010000e-07 V_low
+ 9.000000000e-07 V_low
+ 9.000010000e-07 V_low
+ 9.001000000e-07 V_low
+ 9.001010000e-07 V_low
+ 9.002000000e-07 V_low
+ 9.002010000e-07 V_low
+ 9.003000000e-07 V_low
+ 9.003010000e-07 V_low
+ 9.004000000e-07 V_low
+ 9.004010000e-07 V_low
+ 9.005000000e-07 V_low
+ 9.005010000e-07 V_low
+ 9.006000000e-07 V_low
+ 9.006010000e-07 V_low
+ 9.007000000e-07 V_low
+ 9.007010000e-07 V_low
+ 9.008000000e-07 V_low
+ 9.008010000e-07 V_low
+ 9.009000000e-07 V_low
+ 9.009010000e-07 V_hig
+ 9.010000000e-07 V_hig
+ 9.010010000e-07 V_hig
+ 9.011000000e-07 V_hig
+ 9.011010000e-07 V_hig
+ 9.012000000e-07 V_hig
+ 9.012010000e-07 V_hig
+ 9.013000000e-07 V_hig
+ 9.013010000e-07 V_hig
+ 9.014000000e-07 V_hig
+ 9.014010000e-07 V_hig
+ 9.015000000e-07 V_hig
+ 9.015010000e-07 V_hig
+ 9.016000000e-07 V_hig
+ 9.016010000e-07 V_hig
+ 9.017000000e-07 V_hig
+ 9.017010000e-07 V_hig
+ 9.018000000e-07 V_hig
+ 9.018010000e-07 V_hig
+ 9.019000000e-07 V_hig
+ 9.019010000e-07 V_hig
+ 9.020000000e-07 V_hig
+ 9.020010000e-07 V_hig
+ 9.021000000e-07 V_hig
+ 9.021010000e-07 V_hig
+ 9.022000000e-07 V_hig
+ 9.022010000e-07 V_hig
+ 9.023000000e-07 V_hig
+ 9.023010000e-07 V_hig
+ 9.024000000e-07 V_hig
+ 9.024010000e-07 V_hig
+ 9.025000000e-07 V_hig
+ 9.025010000e-07 V_hig
+ 9.026000000e-07 V_hig
+ 9.026010000e-07 V_hig
+ 9.027000000e-07 V_hig
+ 9.027010000e-07 V_hig
+ 9.028000000e-07 V_hig
+ 9.028010000e-07 V_hig
+ 9.029000000e-07 V_hig
+ 9.029010000e-07 V_hig
+ 9.030000000e-07 V_hig
+ 9.030010000e-07 V_hig
+ 9.031000000e-07 V_hig
+ 9.031010000e-07 V_hig
+ 9.032000000e-07 V_hig
+ 9.032010000e-07 V_hig
+ 9.033000000e-07 V_hig
+ 9.033010000e-07 V_hig
+ 9.034000000e-07 V_hig
+ 9.034010000e-07 V_hig
+ 9.035000000e-07 V_hig
+ 9.035010000e-07 V_hig
+ 9.036000000e-07 V_hig
+ 9.036010000e-07 V_hig
+ 9.037000000e-07 V_hig
+ 9.037010000e-07 V_hig
+ 9.038000000e-07 V_hig
+ 9.038010000e-07 V_hig
+ 9.039000000e-07 V_hig
+ 9.039010000e-07 V_low
+ 9.040000000e-07 V_low
+ 9.040010000e-07 V_low
+ 9.041000000e-07 V_low
+ 9.041010000e-07 V_low
+ 9.042000000e-07 V_low
+ 9.042010000e-07 V_low
+ 9.043000000e-07 V_low
+ 9.043010000e-07 V_low
+ 9.044000000e-07 V_low
+ 9.044010000e-07 V_low
+ 9.045000000e-07 V_low
+ 9.045010000e-07 V_low
+ 9.046000000e-07 V_low
+ 9.046010000e-07 V_low
+ 9.047000000e-07 V_low
+ 9.047010000e-07 V_low
+ 9.048000000e-07 V_low
+ 9.048010000e-07 V_low
+ 9.049000000e-07 V_low
+ 9.049010000e-07 V_low
+ 9.050000000e-07 V_low
+ 9.050010000e-07 V_low
+ 9.051000000e-07 V_low
+ 9.051010000e-07 V_low
+ 9.052000000e-07 V_low
+ 9.052010000e-07 V_low
+ 9.053000000e-07 V_low
+ 9.053010000e-07 V_low
+ 9.054000000e-07 V_low
+ 9.054010000e-07 V_low
+ 9.055000000e-07 V_low
+ 9.055010000e-07 V_low
+ 9.056000000e-07 V_low
+ 9.056010000e-07 V_low
+ 9.057000000e-07 V_low
+ 9.057010000e-07 V_low
+ 9.058000000e-07 V_low
+ 9.058010000e-07 V_low
+ 9.059000000e-07 V_low
+ 9.059010000e-07 V_low
+ 9.060000000e-07 V_low
+ 9.060010000e-07 V_low
+ 9.061000000e-07 V_low
+ 9.061010000e-07 V_low
+ 9.062000000e-07 V_low
+ 9.062010000e-07 V_low
+ 9.063000000e-07 V_low
+ 9.063010000e-07 V_low
+ 9.064000000e-07 V_low
+ 9.064010000e-07 V_low
+ 9.065000000e-07 V_low
+ 9.065010000e-07 V_low
+ 9.066000000e-07 V_low
+ 9.066010000e-07 V_low
+ 9.067000000e-07 V_low
+ 9.067010000e-07 V_low
+ 9.068000000e-07 V_low
+ 9.068010000e-07 V_low
+ 9.069000000e-07 V_low
+ 9.069010000e-07 V_hig
+ 9.070000000e-07 V_hig
+ 9.070010000e-07 V_hig
+ 9.071000000e-07 V_hig
+ 9.071010000e-07 V_hig
+ 9.072000000e-07 V_hig
+ 9.072010000e-07 V_hig
+ 9.073000000e-07 V_hig
+ 9.073010000e-07 V_hig
+ 9.074000000e-07 V_hig
+ 9.074010000e-07 V_hig
+ 9.075000000e-07 V_hig
+ 9.075010000e-07 V_hig
+ 9.076000000e-07 V_hig
+ 9.076010000e-07 V_hig
+ 9.077000000e-07 V_hig
+ 9.077010000e-07 V_hig
+ 9.078000000e-07 V_hig
+ 9.078010000e-07 V_hig
+ 9.079000000e-07 V_hig
+ 9.079010000e-07 V_hig
+ 9.080000000e-07 V_hig
+ 9.080010000e-07 V_hig
+ 9.081000000e-07 V_hig
+ 9.081010000e-07 V_hig
+ 9.082000000e-07 V_hig
+ 9.082010000e-07 V_hig
+ 9.083000000e-07 V_hig
+ 9.083010000e-07 V_hig
+ 9.084000000e-07 V_hig
+ 9.084010000e-07 V_hig
+ 9.085000000e-07 V_hig
+ 9.085010000e-07 V_hig
+ 9.086000000e-07 V_hig
+ 9.086010000e-07 V_hig
+ 9.087000000e-07 V_hig
+ 9.087010000e-07 V_hig
+ 9.088000000e-07 V_hig
+ 9.088010000e-07 V_hig
+ 9.089000000e-07 V_hig
+ 9.089010000e-07 V_low
+ 9.090000000e-07 V_low
+ 9.090010000e-07 V_low
+ 9.091000000e-07 V_low
+ 9.091010000e-07 V_low
+ 9.092000000e-07 V_low
+ 9.092010000e-07 V_low
+ 9.093000000e-07 V_low
+ 9.093010000e-07 V_low
+ 9.094000000e-07 V_low
+ 9.094010000e-07 V_low
+ 9.095000000e-07 V_low
+ 9.095010000e-07 V_low
+ 9.096000000e-07 V_low
+ 9.096010000e-07 V_low
+ 9.097000000e-07 V_low
+ 9.097010000e-07 V_low
+ 9.098000000e-07 V_low
+ 9.098010000e-07 V_low
+ 9.099000000e-07 V_low
+ 9.099010000e-07 V_low
+ 9.100000000e-07 V_low
+ 9.100010000e-07 V_low
+ 9.101000000e-07 V_low
+ 9.101010000e-07 V_low
+ 9.102000000e-07 V_low
+ 9.102010000e-07 V_low
+ 9.103000000e-07 V_low
+ 9.103010000e-07 V_low
+ 9.104000000e-07 V_low
+ 9.104010000e-07 V_low
+ 9.105000000e-07 V_low
+ 9.105010000e-07 V_low
+ 9.106000000e-07 V_low
+ 9.106010000e-07 V_low
+ 9.107000000e-07 V_low
+ 9.107010000e-07 V_low
+ 9.108000000e-07 V_low
+ 9.108010000e-07 V_low
+ 9.109000000e-07 V_low
+ 9.109010000e-07 V_hig
+ 9.110000000e-07 V_hig
+ 9.110010000e-07 V_hig
+ 9.111000000e-07 V_hig
+ 9.111010000e-07 V_hig
+ 9.112000000e-07 V_hig
+ 9.112010000e-07 V_hig
+ 9.113000000e-07 V_hig
+ 9.113010000e-07 V_hig
+ 9.114000000e-07 V_hig
+ 9.114010000e-07 V_hig
+ 9.115000000e-07 V_hig
+ 9.115010000e-07 V_hig
+ 9.116000000e-07 V_hig
+ 9.116010000e-07 V_hig
+ 9.117000000e-07 V_hig
+ 9.117010000e-07 V_hig
+ 9.118000000e-07 V_hig
+ 9.118010000e-07 V_hig
+ 9.119000000e-07 V_hig
+ 9.119010000e-07 V_low
+ 9.120000000e-07 V_low
+ 9.120010000e-07 V_low
+ 9.121000000e-07 V_low
+ 9.121010000e-07 V_low
+ 9.122000000e-07 V_low
+ 9.122010000e-07 V_low
+ 9.123000000e-07 V_low
+ 9.123010000e-07 V_low
+ 9.124000000e-07 V_low
+ 9.124010000e-07 V_low
+ 9.125000000e-07 V_low
+ 9.125010000e-07 V_low
+ 9.126000000e-07 V_low
+ 9.126010000e-07 V_low
+ 9.127000000e-07 V_low
+ 9.127010000e-07 V_low
+ 9.128000000e-07 V_low
+ 9.128010000e-07 V_low
+ 9.129000000e-07 V_low
+ 9.129010000e-07 V_low
+ 9.130000000e-07 V_low
+ 9.130010000e-07 V_low
+ 9.131000000e-07 V_low
+ 9.131010000e-07 V_low
+ 9.132000000e-07 V_low
+ 9.132010000e-07 V_low
+ 9.133000000e-07 V_low
+ 9.133010000e-07 V_low
+ 9.134000000e-07 V_low
+ 9.134010000e-07 V_low
+ 9.135000000e-07 V_low
+ 9.135010000e-07 V_low
+ 9.136000000e-07 V_low
+ 9.136010000e-07 V_low
+ 9.137000000e-07 V_low
+ 9.137010000e-07 V_low
+ 9.138000000e-07 V_low
+ 9.138010000e-07 V_low
+ 9.139000000e-07 V_low
+ 9.139010000e-07 V_low
+ 9.140000000e-07 V_low
+ 9.140010000e-07 V_low
+ 9.141000000e-07 V_low
+ 9.141010000e-07 V_low
+ 9.142000000e-07 V_low
+ 9.142010000e-07 V_low
+ 9.143000000e-07 V_low
+ 9.143010000e-07 V_low
+ 9.144000000e-07 V_low
+ 9.144010000e-07 V_low
+ 9.145000000e-07 V_low
+ 9.145010000e-07 V_low
+ 9.146000000e-07 V_low
+ 9.146010000e-07 V_low
+ 9.147000000e-07 V_low
+ 9.147010000e-07 V_low
+ 9.148000000e-07 V_low
+ 9.148010000e-07 V_low
+ 9.149000000e-07 V_low
+ 9.149010000e-07 V_hig
+ 9.150000000e-07 V_hig
+ 9.150010000e-07 V_hig
+ 9.151000000e-07 V_hig
+ 9.151010000e-07 V_hig
+ 9.152000000e-07 V_hig
+ 9.152010000e-07 V_hig
+ 9.153000000e-07 V_hig
+ 9.153010000e-07 V_hig
+ 9.154000000e-07 V_hig
+ 9.154010000e-07 V_hig
+ 9.155000000e-07 V_hig
+ 9.155010000e-07 V_hig
+ 9.156000000e-07 V_hig
+ 9.156010000e-07 V_hig
+ 9.157000000e-07 V_hig
+ 9.157010000e-07 V_hig
+ 9.158000000e-07 V_hig
+ 9.158010000e-07 V_hig
+ 9.159000000e-07 V_hig
+ 9.159010000e-07 V_hig
+ 9.160000000e-07 V_hig
+ 9.160010000e-07 V_hig
+ 9.161000000e-07 V_hig
+ 9.161010000e-07 V_hig
+ 9.162000000e-07 V_hig
+ 9.162010000e-07 V_hig
+ 9.163000000e-07 V_hig
+ 9.163010000e-07 V_hig
+ 9.164000000e-07 V_hig
+ 9.164010000e-07 V_hig
+ 9.165000000e-07 V_hig
+ 9.165010000e-07 V_hig
+ 9.166000000e-07 V_hig
+ 9.166010000e-07 V_hig
+ 9.167000000e-07 V_hig
+ 9.167010000e-07 V_hig
+ 9.168000000e-07 V_hig
+ 9.168010000e-07 V_hig
+ 9.169000000e-07 V_hig
+ 9.169010000e-07 V_hig
+ 9.170000000e-07 V_hig
+ 9.170010000e-07 V_hig
+ 9.171000000e-07 V_hig
+ 9.171010000e-07 V_hig
+ 9.172000000e-07 V_hig
+ 9.172010000e-07 V_hig
+ 9.173000000e-07 V_hig
+ 9.173010000e-07 V_hig
+ 9.174000000e-07 V_hig
+ 9.174010000e-07 V_hig
+ 9.175000000e-07 V_hig
+ 9.175010000e-07 V_hig
+ 9.176000000e-07 V_hig
+ 9.176010000e-07 V_hig
+ 9.177000000e-07 V_hig
+ 9.177010000e-07 V_hig
+ 9.178000000e-07 V_hig
+ 9.178010000e-07 V_hig
+ 9.179000000e-07 V_hig
+ 9.179010000e-07 V_low
+ 9.180000000e-07 V_low
+ 9.180010000e-07 V_low
+ 9.181000000e-07 V_low
+ 9.181010000e-07 V_low
+ 9.182000000e-07 V_low
+ 9.182010000e-07 V_low
+ 9.183000000e-07 V_low
+ 9.183010000e-07 V_low
+ 9.184000000e-07 V_low
+ 9.184010000e-07 V_low
+ 9.185000000e-07 V_low
+ 9.185010000e-07 V_low
+ 9.186000000e-07 V_low
+ 9.186010000e-07 V_low
+ 9.187000000e-07 V_low
+ 9.187010000e-07 V_low
+ 9.188000000e-07 V_low
+ 9.188010000e-07 V_low
+ 9.189000000e-07 V_low
+ 9.189010000e-07 V_hig
+ 9.190000000e-07 V_hig
+ 9.190010000e-07 V_hig
+ 9.191000000e-07 V_hig
+ 9.191010000e-07 V_hig
+ 9.192000000e-07 V_hig
+ 9.192010000e-07 V_hig
+ 9.193000000e-07 V_hig
+ 9.193010000e-07 V_hig
+ 9.194000000e-07 V_hig
+ 9.194010000e-07 V_hig
+ 9.195000000e-07 V_hig
+ 9.195010000e-07 V_hig
+ 9.196000000e-07 V_hig
+ 9.196010000e-07 V_hig
+ 9.197000000e-07 V_hig
+ 9.197010000e-07 V_hig
+ 9.198000000e-07 V_hig
+ 9.198010000e-07 V_hig
+ 9.199000000e-07 V_hig
+ 9.199010000e-07 V_low
+ 9.200000000e-07 V_low
+ 9.200010000e-07 V_low
+ 9.201000000e-07 V_low
+ 9.201010000e-07 V_low
+ 9.202000000e-07 V_low
+ 9.202010000e-07 V_low
+ 9.203000000e-07 V_low
+ 9.203010000e-07 V_low
+ 9.204000000e-07 V_low
+ 9.204010000e-07 V_low
+ 9.205000000e-07 V_low
+ 9.205010000e-07 V_low
+ 9.206000000e-07 V_low
+ 9.206010000e-07 V_low
+ 9.207000000e-07 V_low
+ 9.207010000e-07 V_low
+ 9.208000000e-07 V_low
+ 9.208010000e-07 V_low
+ 9.209000000e-07 V_low
+ 9.209010000e-07 V_low
+ 9.210000000e-07 V_low
+ 9.210010000e-07 V_low
+ 9.211000000e-07 V_low
+ 9.211010000e-07 V_low
+ 9.212000000e-07 V_low
+ 9.212010000e-07 V_low
+ 9.213000000e-07 V_low
+ 9.213010000e-07 V_low
+ 9.214000000e-07 V_low
+ 9.214010000e-07 V_low
+ 9.215000000e-07 V_low
+ 9.215010000e-07 V_low
+ 9.216000000e-07 V_low
+ 9.216010000e-07 V_low
+ 9.217000000e-07 V_low
+ 9.217010000e-07 V_low
+ 9.218000000e-07 V_low
+ 9.218010000e-07 V_low
+ 9.219000000e-07 V_low
+ 9.219010000e-07 V_low
+ 9.220000000e-07 V_low
+ 9.220010000e-07 V_low
+ 9.221000000e-07 V_low
+ 9.221010000e-07 V_low
+ 9.222000000e-07 V_low
+ 9.222010000e-07 V_low
+ 9.223000000e-07 V_low
+ 9.223010000e-07 V_low
+ 9.224000000e-07 V_low
+ 9.224010000e-07 V_low
+ 9.225000000e-07 V_low
+ 9.225010000e-07 V_low
+ 9.226000000e-07 V_low
+ 9.226010000e-07 V_low
+ 9.227000000e-07 V_low
+ 9.227010000e-07 V_low
+ 9.228000000e-07 V_low
+ 9.228010000e-07 V_low
+ 9.229000000e-07 V_low
+ 9.229010000e-07 V_hig
+ 9.230000000e-07 V_hig
+ 9.230010000e-07 V_hig
+ 9.231000000e-07 V_hig
+ 9.231010000e-07 V_hig
+ 9.232000000e-07 V_hig
+ 9.232010000e-07 V_hig
+ 9.233000000e-07 V_hig
+ 9.233010000e-07 V_hig
+ 9.234000000e-07 V_hig
+ 9.234010000e-07 V_hig
+ 9.235000000e-07 V_hig
+ 9.235010000e-07 V_hig
+ 9.236000000e-07 V_hig
+ 9.236010000e-07 V_hig
+ 9.237000000e-07 V_hig
+ 9.237010000e-07 V_hig
+ 9.238000000e-07 V_hig
+ 9.238010000e-07 V_hig
+ 9.239000000e-07 V_hig
+ 9.239010000e-07 V_low
+ 9.240000000e-07 V_low
+ 9.240010000e-07 V_low
+ 9.241000000e-07 V_low
+ 9.241010000e-07 V_low
+ 9.242000000e-07 V_low
+ 9.242010000e-07 V_low
+ 9.243000000e-07 V_low
+ 9.243010000e-07 V_low
+ 9.244000000e-07 V_low
+ 9.244010000e-07 V_low
+ 9.245000000e-07 V_low
+ 9.245010000e-07 V_low
+ 9.246000000e-07 V_low
+ 9.246010000e-07 V_low
+ 9.247000000e-07 V_low
+ 9.247010000e-07 V_low
+ 9.248000000e-07 V_low
+ 9.248010000e-07 V_low
+ 9.249000000e-07 V_low
+ 9.249010000e-07 V_low
+ 9.250000000e-07 V_low
+ 9.250010000e-07 V_low
+ 9.251000000e-07 V_low
+ 9.251010000e-07 V_low
+ 9.252000000e-07 V_low
+ 9.252010000e-07 V_low
+ 9.253000000e-07 V_low
+ 9.253010000e-07 V_low
+ 9.254000000e-07 V_low
+ 9.254010000e-07 V_low
+ 9.255000000e-07 V_low
+ 9.255010000e-07 V_low
+ 9.256000000e-07 V_low
+ 9.256010000e-07 V_low
+ 9.257000000e-07 V_low
+ 9.257010000e-07 V_low
+ 9.258000000e-07 V_low
+ 9.258010000e-07 V_low
+ 9.259000000e-07 V_low
+ 9.259010000e-07 V_low
+ 9.260000000e-07 V_low
+ 9.260010000e-07 V_low
+ 9.261000000e-07 V_low
+ 9.261010000e-07 V_low
+ 9.262000000e-07 V_low
+ 9.262010000e-07 V_low
+ 9.263000000e-07 V_low
+ 9.263010000e-07 V_low
+ 9.264000000e-07 V_low
+ 9.264010000e-07 V_low
+ 9.265000000e-07 V_low
+ 9.265010000e-07 V_low
+ 9.266000000e-07 V_low
+ 9.266010000e-07 V_low
+ 9.267000000e-07 V_low
+ 9.267010000e-07 V_low
+ 9.268000000e-07 V_low
+ 9.268010000e-07 V_low
+ 9.269000000e-07 V_low
+ 9.269010000e-07 V_hig
+ 9.270000000e-07 V_hig
+ 9.270010000e-07 V_hig
+ 9.271000000e-07 V_hig
+ 9.271010000e-07 V_hig
+ 9.272000000e-07 V_hig
+ 9.272010000e-07 V_hig
+ 9.273000000e-07 V_hig
+ 9.273010000e-07 V_hig
+ 9.274000000e-07 V_hig
+ 9.274010000e-07 V_hig
+ 9.275000000e-07 V_hig
+ 9.275010000e-07 V_hig
+ 9.276000000e-07 V_hig
+ 9.276010000e-07 V_hig
+ 9.277000000e-07 V_hig
+ 9.277010000e-07 V_hig
+ 9.278000000e-07 V_hig
+ 9.278010000e-07 V_hig
+ 9.279000000e-07 V_hig
+ 9.279010000e-07 V_hig
+ 9.280000000e-07 V_hig
+ 9.280010000e-07 V_hig
+ 9.281000000e-07 V_hig
+ 9.281010000e-07 V_hig
+ 9.282000000e-07 V_hig
+ 9.282010000e-07 V_hig
+ 9.283000000e-07 V_hig
+ 9.283010000e-07 V_hig
+ 9.284000000e-07 V_hig
+ 9.284010000e-07 V_hig
+ 9.285000000e-07 V_hig
+ 9.285010000e-07 V_hig
+ 9.286000000e-07 V_hig
+ 9.286010000e-07 V_hig
+ 9.287000000e-07 V_hig
+ 9.287010000e-07 V_hig
+ 9.288000000e-07 V_hig
+ 9.288010000e-07 V_hig
+ 9.289000000e-07 V_hig
+ 9.289010000e-07 V_hig
+ 9.290000000e-07 V_hig
+ 9.290010000e-07 V_hig
+ 9.291000000e-07 V_hig
+ 9.291010000e-07 V_hig
+ 9.292000000e-07 V_hig
+ 9.292010000e-07 V_hig
+ 9.293000000e-07 V_hig
+ 9.293010000e-07 V_hig
+ 9.294000000e-07 V_hig
+ 9.294010000e-07 V_hig
+ 9.295000000e-07 V_hig
+ 9.295010000e-07 V_hig
+ 9.296000000e-07 V_hig
+ 9.296010000e-07 V_hig
+ 9.297000000e-07 V_hig
+ 9.297010000e-07 V_hig
+ 9.298000000e-07 V_hig
+ 9.298010000e-07 V_hig
+ 9.299000000e-07 V_hig
+ 9.299010000e-07 V_hig
+ 9.300000000e-07 V_hig
+ 9.300010000e-07 V_hig
+ 9.301000000e-07 V_hig
+ 9.301010000e-07 V_hig
+ 9.302000000e-07 V_hig
+ 9.302010000e-07 V_hig
+ 9.303000000e-07 V_hig
+ 9.303010000e-07 V_hig
+ 9.304000000e-07 V_hig
+ 9.304010000e-07 V_hig
+ 9.305000000e-07 V_hig
+ 9.305010000e-07 V_hig
+ 9.306000000e-07 V_hig
+ 9.306010000e-07 V_hig
+ 9.307000000e-07 V_hig
+ 9.307010000e-07 V_hig
+ 9.308000000e-07 V_hig
+ 9.308010000e-07 V_hig
+ 9.309000000e-07 V_hig
+ 9.309010000e-07 V_hig
+ 9.310000000e-07 V_hig
+ 9.310010000e-07 V_hig
+ 9.311000000e-07 V_hig
+ 9.311010000e-07 V_hig
+ 9.312000000e-07 V_hig
+ 9.312010000e-07 V_hig
+ 9.313000000e-07 V_hig
+ 9.313010000e-07 V_hig
+ 9.314000000e-07 V_hig
+ 9.314010000e-07 V_hig
+ 9.315000000e-07 V_hig
+ 9.315010000e-07 V_hig
+ 9.316000000e-07 V_hig
+ 9.316010000e-07 V_hig
+ 9.317000000e-07 V_hig
+ 9.317010000e-07 V_hig
+ 9.318000000e-07 V_hig
+ 9.318010000e-07 V_hig
+ 9.319000000e-07 V_hig
+ 9.319010000e-07 V_low
+ 9.320000000e-07 V_low
+ 9.320010000e-07 V_low
+ 9.321000000e-07 V_low
+ 9.321010000e-07 V_low
+ 9.322000000e-07 V_low
+ 9.322010000e-07 V_low
+ 9.323000000e-07 V_low
+ 9.323010000e-07 V_low
+ 9.324000000e-07 V_low
+ 9.324010000e-07 V_low
+ 9.325000000e-07 V_low
+ 9.325010000e-07 V_low
+ 9.326000000e-07 V_low
+ 9.326010000e-07 V_low
+ 9.327000000e-07 V_low
+ 9.327010000e-07 V_low
+ 9.328000000e-07 V_low
+ 9.328010000e-07 V_low
+ 9.329000000e-07 V_low
+ 9.329010000e-07 V_low
+ 9.330000000e-07 V_low
+ 9.330010000e-07 V_low
+ 9.331000000e-07 V_low
+ 9.331010000e-07 V_low
+ 9.332000000e-07 V_low
+ 9.332010000e-07 V_low
+ 9.333000000e-07 V_low
+ 9.333010000e-07 V_low
+ 9.334000000e-07 V_low
+ 9.334010000e-07 V_low
+ 9.335000000e-07 V_low
+ 9.335010000e-07 V_low
+ 9.336000000e-07 V_low
+ 9.336010000e-07 V_low
+ 9.337000000e-07 V_low
+ 9.337010000e-07 V_low
+ 9.338000000e-07 V_low
+ 9.338010000e-07 V_low
+ 9.339000000e-07 V_low
+ 9.339010000e-07 V_low
+ 9.340000000e-07 V_low
+ 9.340010000e-07 V_low
+ 9.341000000e-07 V_low
+ 9.341010000e-07 V_low
+ 9.342000000e-07 V_low
+ 9.342010000e-07 V_low
+ 9.343000000e-07 V_low
+ 9.343010000e-07 V_low
+ 9.344000000e-07 V_low
+ 9.344010000e-07 V_low
+ 9.345000000e-07 V_low
+ 9.345010000e-07 V_low
+ 9.346000000e-07 V_low
+ 9.346010000e-07 V_low
+ 9.347000000e-07 V_low
+ 9.347010000e-07 V_low
+ 9.348000000e-07 V_low
+ 9.348010000e-07 V_low
+ 9.349000000e-07 V_low
+ 9.349010000e-07 V_low
+ 9.350000000e-07 V_low
+ 9.350010000e-07 V_low
+ 9.351000000e-07 V_low
+ 9.351010000e-07 V_low
+ 9.352000000e-07 V_low
+ 9.352010000e-07 V_low
+ 9.353000000e-07 V_low
+ 9.353010000e-07 V_low
+ 9.354000000e-07 V_low
+ 9.354010000e-07 V_low
+ 9.355000000e-07 V_low
+ 9.355010000e-07 V_low
+ 9.356000000e-07 V_low
+ 9.356010000e-07 V_low
+ 9.357000000e-07 V_low
+ 9.357010000e-07 V_low
+ 9.358000000e-07 V_low
+ 9.358010000e-07 V_low
+ 9.359000000e-07 V_low
+ 9.359010000e-07 V_hig
+ 9.360000000e-07 V_hig
+ 9.360010000e-07 V_hig
+ 9.361000000e-07 V_hig
+ 9.361010000e-07 V_hig
+ 9.362000000e-07 V_hig
+ 9.362010000e-07 V_hig
+ 9.363000000e-07 V_hig
+ 9.363010000e-07 V_hig
+ 9.364000000e-07 V_hig
+ 9.364010000e-07 V_hig
+ 9.365000000e-07 V_hig
+ 9.365010000e-07 V_hig
+ 9.366000000e-07 V_hig
+ 9.366010000e-07 V_hig
+ 9.367000000e-07 V_hig
+ 9.367010000e-07 V_hig
+ 9.368000000e-07 V_hig
+ 9.368010000e-07 V_hig
+ 9.369000000e-07 V_hig
+ 9.369010000e-07 V_hig
+ 9.370000000e-07 V_hig
+ 9.370010000e-07 V_hig
+ 9.371000000e-07 V_hig
+ 9.371010000e-07 V_hig
+ 9.372000000e-07 V_hig
+ 9.372010000e-07 V_hig
+ 9.373000000e-07 V_hig
+ 9.373010000e-07 V_hig
+ 9.374000000e-07 V_hig
+ 9.374010000e-07 V_hig
+ 9.375000000e-07 V_hig
+ 9.375010000e-07 V_hig
+ 9.376000000e-07 V_hig
+ 9.376010000e-07 V_hig
+ 9.377000000e-07 V_hig
+ 9.377010000e-07 V_hig
+ 9.378000000e-07 V_hig
+ 9.378010000e-07 V_hig
+ 9.379000000e-07 V_hig
+ 9.379010000e-07 V_low
+ 9.380000000e-07 V_low
+ 9.380010000e-07 V_low
+ 9.381000000e-07 V_low
+ 9.381010000e-07 V_low
+ 9.382000000e-07 V_low
+ 9.382010000e-07 V_low
+ 9.383000000e-07 V_low
+ 9.383010000e-07 V_low
+ 9.384000000e-07 V_low
+ 9.384010000e-07 V_low
+ 9.385000000e-07 V_low
+ 9.385010000e-07 V_low
+ 9.386000000e-07 V_low
+ 9.386010000e-07 V_low
+ 9.387000000e-07 V_low
+ 9.387010000e-07 V_low
+ 9.388000000e-07 V_low
+ 9.388010000e-07 V_low
+ 9.389000000e-07 V_low
+ 9.389010000e-07 V_low
+ 9.390000000e-07 V_low
+ 9.390010000e-07 V_low
+ 9.391000000e-07 V_low
+ 9.391010000e-07 V_low
+ 9.392000000e-07 V_low
+ 9.392010000e-07 V_low
+ 9.393000000e-07 V_low
+ 9.393010000e-07 V_low
+ 9.394000000e-07 V_low
+ 9.394010000e-07 V_low
+ 9.395000000e-07 V_low
+ 9.395010000e-07 V_low
+ 9.396000000e-07 V_low
+ 9.396010000e-07 V_low
+ 9.397000000e-07 V_low
+ 9.397010000e-07 V_low
+ 9.398000000e-07 V_low
+ 9.398010000e-07 V_low
+ 9.399000000e-07 V_low
+ 9.399010000e-07 V_hig
+ 9.400000000e-07 V_hig
+ 9.400010000e-07 V_hig
+ 9.401000000e-07 V_hig
+ 9.401010000e-07 V_hig
+ 9.402000000e-07 V_hig
+ 9.402010000e-07 V_hig
+ 9.403000000e-07 V_hig
+ 9.403010000e-07 V_hig
+ 9.404000000e-07 V_hig
+ 9.404010000e-07 V_hig
+ 9.405000000e-07 V_hig
+ 9.405010000e-07 V_hig
+ 9.406000000e-07 V_hig
+ 9.406010000e-07 V_hig
+ 9.407000000e-07 V_hig
+ 9.407010000e-07 V_hig
+ 9.408000000e-07 V_hig
+ 9.408010000e-07 V_hig
+ 9.409000000e-07 V_hig
+ 9.409010000e-07 V_hig
+ 9.410000000e-07 V_hig
+ 9.410010000e-07 V_hig
+ 9.411000000e-07 V_hig
+ 9.411010000e-07 V_hig
+ 9.412000000e-07 V_hig
+ 9.412010000e-07 V_hig
+ 9.413000000e-07 V_hig
+ 9.413010000e-07 V_hig
+ 9.414000000e-07 V_hig
+ 9.414010000e-07 V_hig
+ 9.415000000e-07 V_hig
+ 9.415010000e-07 V_hig
+ 9.416000000e-07 V_hig
+ 9.416010000e-07 V_hig
+ 9.417000000e-07 V_hig
+ 9.417010000e-07 V_hig
+ 9.418000000e-07 V_hig
+ 9.418010000e-07 V_hig
+ 9.419000000e-07 V_hig
+ 9.419010000e-07 V_low
+ 9.420000000e-07 V_low
+ 9.420010000e-07 V_low
+ 9.421000000e-07 V_low
+ 9.421010000e-07 V_low
+ 9.422000000e-07 V_low
+ 9.422010000e-07 V_low
+ 9.423000000e-07 V_low
+ 9.423010000e-07 V_low
+ 9.424000000e-07 V_low
+ 9.424010000e-07 V_low
+ 9.425000000e-07 V_low
+ 9.425010000e-07 V_low
+ 9.426000000e-07 V_low
+ 9.426010000e-07 V_low
+ 9.427000000e-07 V_low
+ 9.427010000e-07 V_low
+ 9.428000000e-07 V_low
+ 9.428010000e-07 V_low
+ 9.429000000e-07 V_low
+ 9.429010000e-07 V_low
+ 9.430000000e-07 V_low
+ 9.430010000e-07 V_low
+ 9.431000000e-07 V_low
+ 9.431010000e-07 V_low
+ 9.432000000e-07 V_low
+ 9.432010000e-07 V_low
+ 9.433000000e-07 V_low
+ 9.433010000e-07 V_low
+ 9.434000000e-07 V_low
+ 9.434010000e-07 V_low
+ 9.435000000e-07 V_low
+ 9.435010000e-07 V_low
+ 9.436000000e-07 V_low
+ 9.436010000e-07 V_low
+ 9.437000000e-07 V_low
+ 9.437010000e-07 V_low
+ 9.438000000e-07 V_low
+ 9.438010000e-07 V_low
+ 9.439000000e-07 V_low
+ 9.439010000e-07 V_hig
+ 9.440000000e-07 V_hig
+ 9.440010000e-07 V_hig
+ 9.441000000e-07 V_hig
+ 9.441010000e-07 V_hig
+ 9.442000000e-07 V_hig
+ 9.442010000e-07 V_hig
+ 9.443000000e-07 V_hig
+ 9.443010000e-07 V_hig
+ 9.444000000e-07 V_hig
+ 9.444010000e-07 V_hig
+ 9.445000000e-07 V_hig
+ 9.445010000e-07 V_hig
+ 9.446000000e-07 V_hig
+ 9.446010000e-07 V_hig
+ 9.447000000e-07 V_hig
+ 9.447010000e-07 V_hig
+ 9.448000000e-07 V_hig
+ 9.448010000e-07 V_hig
+ 9.449000000e-07 V_hig
+ 9.449010000e-07 V_hig
+ 9.450000000e-07 V_hig
+ 9.450010000e-07 V_hig
+ 9.451000000e-07 V_hig
+ 9.451010000e-07 V_hig
+ 9.452000000e-07 V_hig
+ 9.452010000e-07 V_hig
+ 9.453000000e-07 V_hig
+ 9.453010000e-07 V_hig
+ 9.454000000e-07 V_hig
+ 9.454010000e-07 V_hig
+ 9.455000000e-07 V_hig
+ 9.455010000e-07 V_hig
+ 9.456000000e-07 V_hig
+ 9.456010000e-07 V_hig
+ 9.457000000e-07 V_hig
+ 9.457010000e-07 V_hig
+ 9.458000000e-07 V_hig
+ 9.458010000e-07 V_hig
+ 9.459000000e-07 V_hig
+ 9.459010000e-07 V_low
+ 9.460000000e-07 V_low
+ 9.460010000e-07 V_low
+ 9.461000000e-07 V_low
+ 9.461010000e-07 V_low
+ 9.462000000e-07 V_low
+ 9.462010000e-07 V_low
+ 9.463000000e-07 V_low
+ 9.463010000e-07 V_low
+ 9.464000000e-07 V_low
+ 9.464010000e-07 V_low
+ 9.465000000e-07 V_low
+ 9.465010000e-07 V_low
+ 9.466000000e-07 V_low
+ 9.466010000e-07 V_low
+ 9.467000000e-07 V_low
+ 9.467010000e-07 V_low
+ 9.468000000e-07 V_low
+ 9.468010000e-07 V_low
+ 9.469000000e-07 V_low
+ 9.469010000e-07 V_low
+ 9.470000000e-07 V_low
+ 9.470010000e-07 V_low
+ 9.471000000e-07 V_low
+ 9.471010000e-07 V_low
+ 9.472000000e-07 V_low
+ 9.472010000e-07 V_low
+ 9.473000000e-07 V_low
+ 9.473010000e-07 V_low
+ 9.474000000e-07 V_low
+ 9.474010000e-07 V_low
+ 9.475000000e-07 V_low
+ 9.475010000e-07 V_low
+ 9.476000000e-07 V_low
+ 9.476010000e-07 V_low
+ 9.477000000e-07 V_low
+ 9.477010000e-07 V_low
+ 9.478000000e-07 V_low
+ 9.478010000e-07 V_low
+ 9.479000000e-07 V_low
+ 9.479010000e-07 V_low
+ 9.480000000e-07 V_low
+ 9.480010000e-07 V_low
+ 9.481000000e-07 V_low
+ 9.481010000e-07 V_low
+ 9.482000000e-07 V_low
+ 9.482010000e-07 V_low
+ 9.483000000e-07 V_low
+ 9.483010000e-07 V_low
+ 9.484000000e-07 V_low
+ 9.484010000e-07 V_low
+ 9.485000000e-07 V_low
+ 9.485010000e-07 V_low
+ 9.486000000e-07 V_low
+ 9.486010000e-07 V_low
+ 9.487000000e-07 V_low
+ 9.487010000e-07 V_low
+ 9.488000000e-07 V_low
+ 9.488010000e-07 V_low
+ 9.489000000e-07 V_low
+ 9.489010000e-07 V_hig
+ 9.490000000e-07 V_hig
+ 9.490010000e-07 V_hig
+ 9.491000000e-07 V_hig
+ 9.491010000e-07 V_hig
+ 9.492000000e-07 V_hig
+ 9.492010000e-07 V_hig
+ 9.493000000e-07 V_hig
+ 9.493010000e-07 V_hig
+ 9.494000000e-07 V_hig
+ 9.494010000e-07 V_hig
+ 9.495000000e-07 V_hig
+ 9.495010000e-07 V_hig
+ 9.496000000e-07 V_hig
+ 9.496010000e-07 V_hig
+ 9.497000000e-07 V_hig
+ 9.497010000e-07 V_hig
+ 9.498000000e-07 V_hig
+ 9.498010000e-07 V_hig
+ 9.499000000e-07 V_hig
+ 9.499010000e-07 V_hig
+ 9.500000000e-07 V_hig
+ 9.500010000e-07 V_hig
+ 9.501000000e-07 V_hig
+ 9.501010000e-07 V_hig
+ 9.502000000e-07 V_hig
+ 9.502010000e-07 V_hig
+ 9.503000000e-07 V_hig
+ 9.503010000e-07 V_hig
+ 9.504000000e-07 V_hig
+ 9.504010000e-07 V_hig
+ 9.505000000e-07 V_hig
+ 9.505010000e-07 V_hig
+ 9.506000000e-07 V_hig
+ 9.506010000e-07 V_hig
+ 9.507000000e-07 V_hig
+ 9.507010000e-07 V_hig
+ 9.508000000e-07 V_hig
+ 9.508010000e-07 V_hig
+ 9.509000000e-07 V_hig
+ 9.509010000e-07 V_low
+ 9.510000000e-07 V_low
+ 9.510010000e-07 V_low
+ 9.511000000e-07 V_low
+ 9.511010000e-07 V_low
+ 9.512000000e-07 V_low
+ 9.512010000e-07 V_low
+ 9.513000000e-07 V_low
+ 9.513010000e-07 V_low
+ 9.514000000e-07 V_low
+ 9.514010000e-07 V_low
+ 9.515000000e-07 V_low
+ 9.515010000e-07 V_low
+ 9.516000000e-07 V_low
+ 9.516010000e-07 V_low
+ 9.517000000e-07 V_low
+ 9.517010000e-07 V_low
+ 9.518000000e-07 V_low
+ 9.518010000e-07 V_low
+ 9.519000000e-07 V_low
+ 9.519010000e-07 V_low
+ 9.520000000e-07 V_low
+ 9.520010000e-07 V_low
+ 9.521000000e-07 V_low
+ 9.521010000e-07 V_low
+ 9.522000000e-07 V_low
+ 9.522010000e-07 V_low
+ 9.523000000e-07 V_low
+ 9.523010000e-07 V_low
+ 9.524000000e-07 V_low
+ 9.524010000e-07 V_low
+ 9.525000000e-07 V_low
+ 9.525010000e-07 V_low
+ 9.526000000e-07 V_low
+ 9.526010000e-07 V_low
+ 9.527000000e-07 V_low
+ 9.527010000e-07 V_low
+ 9.528000000e-07 V_low
+ 9.528010000e-07 V_low
+ 9.529000000e-07 V_low
+ 9.529010000e-07 V_hig
+ 9.530000000e-07 V_hig
+ 9.530010000e-07 V_hig
+ 9.531000000e-07 V_hig
+ 9.531010000e-07 V_hig
+ 9.532000000e-07 V_hig
+ 9.532010000e-07 V_hig
+ 9.533000000e-07 V_hig
+ 9.533010000e-07 V_hig
+ 9.534000000e-07 V_hig
+ 9.534010000e-07 V_hig
+ 9.535000000e-07 V_hig
+ 9.535010000e-07 V_hig
+ 9.536000000e-07 V_hig
+ 9.536010000e-07 V_hig
+ 9.537000000e-07 V_hig
+ 9.537010000e-07 V_hig
+ 9.538000000e-07 V_hig
+ 9.538010000e-07 V_hig
+ 9.539000000e-07 V_hig
+ 9.539010000e-07 V_hig
+ 9.540000000e-07 V_hig
+ 9.540010000e-07 V_hig
+ 9.541000000e-07 V_hig
+ 9.541010000e-07 V_hig
+ 9.542000000e-07 V_hig
+ 9.542010000e-07 V_hig
+ 9.543000000e-07 V_hig
+ 9.543010000e-07 V_hig
+ 9.544000000e-07 V_hig
+ 9.544010000e-07 V_hig
+ 9.545000000e-07 V_hig
+ 9.545010000e-07 V_hig
+ 9.546000000e-07 V_hig
+ 9.546010000e-07 V_hig
+ 9.547000000e-07 V_hig
+ 9.547010000e-07 V_hig
+ 9.548000000e-07 V_hig
+ 9.548010000e-07 V_hig
+ 9.549000000e-07 V_hig
+ 9.549010000e-07 V_hig
+ 9.550000000e-07 V_hig
+ 9.550010000e-07 V_hig
+ 9.551000000e-07 V_hig
+ 9.551010000e-07 V_hig
+ 9.552000000e-07 V_hig
+ 9.552010000e-07 V_hig
+ 9.553000000e-07 V_hig
+ 9.553010000e-07 V_hig
+ 9.554000000e-07 V_hig
+ 9.554010000e-07 V_hig
+ 9.555000000e-07 V_hig
+ 9.555010000e-07 V_hig
+ 9.556000000e-07 V_hig
+ 9.556010000e-07 V_hig
+ 9.557000000e-07 V_hig
+ 9.557010000e-07 V_hig
+ 9.558000000e-07 V_hig
+ 9.558010000e-07 V_hig
+ 9.559000000e-07 V_hig
+ 9.559010000e-07 V_low
+ 9.560000000e-07 V_low
+ 9.560010000e-07 V_low
+ 9.561000000e-07 V_low
+ 9.561010000e-07 V_low
+ 9.562000000e-07 V_low
+ 9.562010000e-07 V_low
+ 9.563000000e-07 V_low
+ 9.563010000e-07 V_low
+ 9.564000000e-07 V_low
+ 9.564010000e-07 V_low
+ 9.565000000e-07 V_low
+ 9.565010000e-07 V_low
+ 9.566000000e-07 V_low
+ 9.566010000e-07 V_low
+ 9.567000000e-07 V_low
+ 9.567010000e-07 V_low
+ 9.568000000e-07 V_low
+ 9.568010000e-07 V_low
+ 9.569000000e-07 V_low
+ 9.569010000e-07 V_hig
+ 9.570000000e-07 V_hig
+ 9.570010000e-07 V_hig
+ 9.571000000e-07 V_hig
+ 9.571010000e-07 V_hig
+ 9.572000000e-07 V_hig
+ 9.572010000e-07 V_hig
+ 9.573000000e-07 V_hig
+ 9.573010000e-07 V_hig
+ 9.574000000e-07 V_hig
+ 9.574010000e-07 V_hig
+ 9.575000000e-07 V_hig
+ 9.575010000e-07 V_hig
+ 9.576000000e-07 V_hig
+ 9.576010000e-07 V_hig
+ 9.577000000e-07 V_hig
+ 9.577010000e-07 V_hig
+ 9.578000000e-07 V_hig
+ 9.578010000e-07 V_hig
+ 9.579000000e-07 V_hig
+ 9.579010000e-07 V_hig
+ 9.580000000e-07 V_hig
+ 9.580010000e-07 V_hig
+ 9.581000000e-07 V_hig
+ 9.581010000e-07 V_hig
+ 9.582000000e-07 V_hig
+ 9.582010000e-07 V_hig
+ 9.583000000e-07 V_hig
+ 9.583010000e-07 V_hig
+ 9.584000000e-07 V_hig
+ 9.584010000e-07 V_hig
+ 9.585000000e-07 V_hig
+ 9.585010000e-07 V_hig
+ 9.586000000e-07 V_hig
+ 9.586010000e-07 V_hig
+ 9.587000000e-07 V_hig
+ 9.587010000e-07 V_hig
+ 9.588000000e-07 V_hig
+ 9.588010000e-07 V_hig
+ 9.589000000e-07 V_hig
+ 9.589010000e-07 V_low
+ 9.590000000e-07 V_low
+ 9.590010000e-07 V_low
+ 9.591000000e-07 V_low
+ 9.591010000e-07 V_low
+ 9.592000000e-07 V_low
+ 9.592010000e-07 V_low
+ 9.593000000e-07 V_low
+ 9.593010000e-07 V_low
+ 9.594000000e-07 V_low
+ 9.594010000e-07 V_low
+ 9.595000000e-07 V_low
+ 9.595010000e-07 V_low
+ 9.596000000e-07 V_low
+ 9.596010000e-07 V_low
+ 9.597000000e-07 V_low
+ 9.597010000e-07 V_low
+ 9.598000000e-07 V_low
+ 9.598010000e-07 V_low
+ 9.599000000e-07 V_low
+ 9.599010000e-07 V_hig
+ 9.600000000e-07 V_hig
+ 9.600010000e-07 V_hig
+ 9.601000000e-07 V_hig
+ 9.601010000e-07 V_hig
+ 9.602000000e-07 V_hig
+ 9.602010000e-07 V_hig
+ 9.603000000e-07 V_hig
+ 9.603010000e-07 V_hig
+ 9.604000000e-07 V_hig
+ 9.604010000e-07 V_hig
+ 9.605000000e-07 V_hig
+ 9.605010000e-07 V_hig
+ 9.606000000e-07 V_hig
+ 9.606010000e-07 V_hig
+ 9.607000000e-07 V_hig
+ 9.607010000e-07 V_hig
+ 9.608000000e-07 V_hig
+ 9.608010000e-07 V_hig
+ 9.609000000e-07 V_hig
+ 9.609010000e-07 V_hig
+ 9.610000000e-07 V_hig
+ 9.610010000e-07 V_hig
+ 9.611000000e-07 V_hig
+ 9.611010000e-07 V_hig
+ 9.612000000e-07 V_hig
+ 9.612010000e-07 V_hig
+ 9.613000000e-07 V_hig
+ 9.613010000e-07 V_hig
+ 9.614000000e-07 V_hig
+ 9.614010000e-07 V_hig
+ 9.615000000e-07 V_hig
+ 9.615010000e-07 V_hig
+ 9.616000000e-07 V_hig
+ 9.616010000e-07 V_hig
+ 9.617000000e-07 V_hig
+ 9.617010000e-07 V_hig
+ 9.618000000e-07 V_hig
+ 9.618010000e-07 V_hig
+ 9.619000000e-07 V_hig
+ 9.619010000e-07 V_hig
+ 9.620000000e-07 V_hig
+ 9.620010000e-07 V_hig
+ 9.621000000e-07 V_hig
+ 9.621010000e-07 V_hig
+ 9.622000000e-07 V_hig
+ 9.622010000e-07 V_hig
+ 9.623000000e-07 V_hig
+ 9.623010000e-07 V_hig
+ 9.624000000e-07 V_hig
+ 9.624010000e-07 V_hig
+ 9.625000000e-07 V_hig
+ 9.625010000e-07 V_hig
+ 9.626000000e-07 V_hig
+ 9.626010000e-07 V_hig
+ 9.627000000e-07 V_hig
+ 9.627010000e-07 V_hig
+ 9.628000000e-07 V_hig
+ 9.628010000e-07 V_hig
+ 9.629000000e-07 V_hig
+ 9.629010000e-07 V_hig
+ 9.630000000e-07 V_hig
+ 9.630010000e-07 V_hig
+ 9.631000000e-07 V_hig
+ 9.631010000e-07 V_hig
+ 9.632000000e-07 V_hig
+ 9.632010000e-07 V_hig
+ 9.633000000e-07 V_hig
+ 9.633010000e-07 V_hig
+ 9.634000000e-07 V_hig
+ 9.634010000e-07 V_hig
+ 9.635000000e-07 V_hig
+ 9.635010000e-07 V_hig
+ 9.636000000e-07 V_hig
+ 9.636010000e-07 V_hig
+ 9.637000000e-07 V_hig
+ 9.637010000e-07 V_hig
+ 9.638000000e-07 V_hig
+ 9.638010000e-07 V_hig
+ 9.639000000e-07 V_hig
+ 9.639010000e-07 V_low
+ 9.640000000e-07 V_low
+ 9.640010000e-07 V_low
+ 9.641000000e-07 V_low
+ 9.641010000e-07 V_low
+ 9.642000000e-07 V_low
+ 9.642010000e-07 V_low
+ 9.643000000e-07 V_low
+ 9.643010000e-07 V_low
+ 9.644000000e-07 V_low
+ 9.644010000e-07 V_low
+ 9.645000000e-07 V_low
+ 9.645010000e-07 V_low
+ 9.646000000e-07 V_low
+ 9.646010000e-07 V_low
+ 9.647000000e-07 V_low
+ 9.647010000e-07 V_low
+ 9.648000000e-07 V_low
+ 9.648010000e-07 V_low
+ 9.649000000e-07 V_low
+ 9.649010000e-07 V_hig
+ 9.650000000e-07 V_hig
+ 9.650010000e-07 V_hig
+ 9.651000000e-07 V_hig
+ 9.651010000e-07 V_hig
+ 9.652000000e-07 V_hig
+ 9.652010000e-07 V_hig
+ 9.653000000e-07 V_hig
+ 9.653010000e-07 V_hig
+ 9.654000000e-07 V_hig
+ 9.654010000e-07 V_hig
+ 9.655000000e-07 V_hig
+ 9.655010000e-07 V_hig
+ 9.656000000e-07 V_hig
+ 9.656010000e-07 V_hig
+ 9.657000000e-07 V_hig
+ 9.657010000e-07 V_hig
+ 9.658000000e-07 V_hig
+ 9.658010000e-07 V_hig
+ 9.659000000e-07 V_hig
+ 9.659010000e-07 V_hig
+ 9.660000000e-07 V_hig
+ 9.660010000e-07 V_hig
+ 9.661000000e-07 V_hig
+ 9.661010000e-07 V_hig
+ 9.662000000e-07 V_hig
+ 9.662010000e-07 V_hig
+ 9.663000000e-07 V_hig
+ 9.663010000e-07 V_hig
+ 9.664000000e-07 V_hig
+ 9.664010000e-07 V_hig
+ 9.665000000e-07 V_hig
+ 9.665010000e-07 V_hig
+ 9.666000000e-07 V_hig
+ 9.666010000e-07 V_hig
+ 9.667000000e-07 V_hig
+ 9.667010000e-07 V_hig
+ 9.668000000e-07 V_hig
+ 9.668010000e-07 V_hig
+ 9.669000000e-07 V_hig
+ 9.669010000e-07 V_hig
+ 9.670000000e-07 V_hig
+ 9.670010000e-07 V_hig
+ 9.671000000e-07 V_hig
+ 9.671010000e-07 V_hig
+ 9.672000000e-07 V_hig
+ 9.672010000e-07 V_hig
+ 9.673000000e-07 V_hig
+ 9.673010000e-07 V_hig
+ 9.674000000e-07 V_hig
+ 9.674010000e-07 V_hig
+ 9.675000000e-07 V_hig
+ 9.675010000e-07 V_hig
+ 9.676000000e-07 V_hig
+ 9.676010000e-07 V_hig
+ 9.677000000e-07 V_hig
+ 9.677010000e-07 V_hig
+ 9.678000000e-07 V_hig
+ 9.678010000e-07 V_hig
+ 9.679000000e-07 V_hig
+ 9.679010000e-07 V_low
+ 9.680000000e-07 V_low
+ 9.680010000e-07 V_low
+ 9.681000000e-07 V_low
+ 9.681010000e-07 V_low
+ 9.682000000e-07 V_low
+ 9.682010000e-07 V_low
+ 9.683000000e-07 V_low
+ 9.683010000e-07 V_low
+ 9.684000000e-07 V_low
+ 9.684010000e-07 V_low
+ 9.685000000e-07 V_low
+ 9.685010000e-07 V_low
+ 9.686000000e-07 V_low
+ 9.686010000e-07 V_low
+ 9.687000000e-07 V_low
+ 9.687010000e-07 V_low
+ 9.688000000e-07 V_low
+ 9.688010000e-07 V_low
+ 9.689000000e-07 V_low
+ 9.689010000e-07 V_low
+ 9.690000000e-07 V_low
+ 9.690010000e-07 V_low
+ 9.691000000e-07 V_low
+ 9.691010000e-07 V_low
+ 9.692000000e-07 V_low
+ 9.692010000e-07 V_low
+ 9.693000000e-07 V_low
+ 9.693010000e-07 V_low
+ 9.694000000e-07 V_low
+ 9.694010000e-07 V_low
+ 9.695000000e-07 V_low
+ 9.695010000e-07 V_low
+ 9.696000000e-07 V_low
+ 9.696010000e-07 V_low
+ 9.697000000e-07 V_low
+ 9.697010000e-07 V_low
+ 9.698000000e-07 V_low
+ 9.698010000e-07 V_low
+ 9.699000000e-07 V_low
+ 9.699010000e-07 V_low
+ 9.700000000e-07 V_low
+ 9.700010000e-07 V_low
+ 9.701000000e-07 V_low
+ 9.701010000e-07 V_low
+ 9.702000000e-07 V_low
+ 9.702010000e-07 V_low
+ 9.703000000e-07 V_low
+ 9.703010000e-07 V_low
+ 9.704000000e-07 V_low
+ 9.704010000e-07 V_low
+ 9.705000000e-07 V_low
+ 9.705010000e-07 V_low
+ 9.706000000e-07 V_low
+ 9.706010000e-07 V_low
+ 9.707000000e-07 V_low
+ 9.707010000e-07 V_low
+ 9.708000000e-07 V_low
+ 9.708010000e-07 V_low
+ 9.709000000e-07 V_low
+ 9.709010000e-07 V_hig
+ 9.710000000e-07 V_hig
+ 9.710010000e-07 V_hig
+ 9.711000000e-07 V_hig
+ 9.711010000e-07 V_hig
+ 9.712000000e-07 V_hig
+ 9.712010000e-07 V_hig
+ 9.713000000e-07 V_hig
+ 9.713010000e-07 V_hig
+ 9.714000000e-07 V_hig
+ 9.714010000e-07 V_hig
+ 9.715000000e-07 V_hig
+ 9.715010000e-07 V_hig
+ 9.716000000e-07 V_hig
+ 9.716010000e-07 V_hig
+ 9.717000000e-07 V_hig
+ 9.717010000e-07 V_hig
+ 9.718000000e-07 V_hig
+ 9.718010000e-07 V_hig
+ 9.719000000e-07 V_hig
+ 9.719010000e-07 V_low
+ 9.720000000e-07 V_low
+ 9.720010000e-07 V_low
+ 9.721000000e-07 V_low
+ 9.721010000e-07 V_low
+ 9.722000000e-07 V_low
+ 9.722010000e-07 V_low
+ 9.723000000e-07 V_low
+ 9.723010000e-07 V_low
+ 9.724000000e-07 V_low
+ 9.724010000e-07 V_low
+ 9.725000000e-07 V_low
+ 9.725010000e-07 V_low
+ 9.726000000e-07 V_low
+ 9.726010000e-07 V_low
+ 9.727000000e-07 V_low
+ 9.727010000e-07 V_low
+ 9.728000000e-07 V_low
+ 9.728010000e-07 V_low
+ 9.729000000e-07 V_low
+ 9.729010000e-07 V_low
+ 9.730000000e-07 V_low
+ 9.730010000e-07 V_low
+ 9.731000000e-07 V_low
+ 9.731010000e-07 V_low
+ 9.732000000e-07 V_low
+ 9.732010000e-07 V_low
+ 9.733000000e-07 V_low
+ 9.733010000e-07 V_low
+ 9.734000000e-07 V_low
+ 9.734010000e-07 V_low
+ 9.735000000e-07 V_low
+ 9.735010000e-07 V_low
+ 9.736000000e-07 V_low
+ 9.736010000e-07 V_low
+ 9.737000000e-07 V_low
+ 9.737010000e-07 V_low
+ 9.738000000e-07 V_low
+ 9.738010000e-07 V_low
+ 9.739000000e-07 V_low
+ 9.739010000e-07 V_low
+ 9.740000000e-07 V_low
+ 9.740010000e-07 V_low
+ 9.741000000e-07 V_low
+ 9.741010000e-07 V_low
+ 9.742000000e-07 V_low
+ 9.742010000e-07 V_low
+ 9.743000000e-07 V_low
+ 9.743010000e-07 V_low
+ 9.744000000e-07 V_low
+ 9.744010000e-07 V_low
+ 9.745000000e-07 V_low
+ 9.745010000e-07 V_low
+ 9.746000000e-07 V_low
+ 9.746010000e-07 V_low
+ 9.747000000e-07 V_low
+ 9.747010000e-07 V_low
+ 9.748000000e-07 V_low
+ 9.748010000e-07 V_low
+ 9.749000000e-07 V_low
+ 9.749010000e-07 V_hig
+ 9.750000000e-07 V_hig
+ 9.750010000e-07 V_hig
+ 9.751000000e-07 V_hig
+ 9.751010000e-07 V_hig
+ 9.752000000e-07 V_hig
+ 9.752010000e-07 V_hig
+ 9.753000000e-07 V_hig
+ 9.753010000e-07 V_hig
+ 9.754000000e-07 V_hig
+ 9.754010000e-07 V_hig
+ 9.755000000e-07 V_hig
+ 9.755010000e-07 V_hig
+ 9.756000000e-07 V_hig
+ 9.756010000e-07 V_hig
+ 9.757000000e-07 V_hig
+ 9.757010000e-07 V_hig
+ 9.758000000e-07 V_hig
+ 9.758010000e-07 V_hig
+ 9.759000000e-07 V_hig
+ 9.759010000e-07 V_hig
+ 9.760000000e-07 V_hig
+ 9.760010000e-07 V_hig
+ 9.761000000e-07 V_hig
+ 9.761010000e-07 V_hig
+ 9.762000000e-07 V_hig
+ 9.762010000e-07 V_hig
+ 9.763000000e-07 V_hig
+ 9.763010000e-07 V_hig
+ 9.764000000e-07 V_hig
+ 9.764010000e-07 V_hig
+ 9.765000000e-07 V_hig
+ 9.765010000e-07 V_hig
+ 9.766000000e-07 V_hig
+ 9.766010000e-07 V_hig
+ 9.767000000e-07 V_hig
+ 9.767010000e-07 V_hig
+ 9.768000000e-07 V_hig
+ 9.768010000e-07 V_hig
+ 9.769000000e-07 V_hig
+ 9.769010000e-07 V_hig
+ 9.770000000e-07 V_hig
+ 9.770010000e-07 V_hig
+ 9.771000000e-07 V_hig
+ 9.771010000e-07 V_hig
+ 9.772000000e-07 V_hig
+ 9.772010000e-07 V_hig
+ 9.773000000e-07 V_hig
+ 9.773010000e-07 V_hig
+ 9.774000000e-07 V_hig
+ 9.774010000e-07 V_hig
+ 9.775000000e-07 V_hig
+ 9.775010000e-07 V_hig
+ 9.776000000e-07 V_hig
+ 9.776010000e-07 V_hig
+ 9.777000000e-07 V_hig
+ 9.777010000e-07 V_hig
+ 9.778000000e-07 V_hig
+ 9.778010000e-07 V_hig
+ 9.779000000e-07 V_hig
+ 9.779010000e-07 V_hig
+ 9.780000000e-07 V_hig
+ 9.780010000e-07 V_hig
+ 9.781000000e-07 V_hig
+ 9.781010000e-07 V_hig
+ 9.782000000e-07 V_hig
+ 9.782010000e-07 V_hig
+ 9.783000000e-07 V_hig
+ 9.783010000e-07 V_hig
+ 9.784000000e-07 V_hig
+ 9.784010000e-07 V_hig
+ 9.785000000e-07 V_hig
+ 9.785010000e-07 V_hig
+ 9.786000000e-07 V_hig
+ 9.786010000e-07 V_hig
+ 9.787000000e-07 V_hig
+ 9.787010000e-07 V_hig
+ 9.788000000e-07 V_hig
+ 9.788010000e-07 V_hig
+ 9.789000000e-07 V_hig
+ 9.789010000e-07 V_low
+ 9.790000000e-07 V_low
+ 9.790010000e-07 V_low
+ 9.791000000e-07 V_low
+ 9.791010000e-07 V_low
+ 9.792000000e-07 V_low
+ 9.792010000e-07 V_low
+ 9.793000000e-07 V_low
+ 9.793010000e-07 V_low
+ 9.794000000e-07 V_low
+ 9.794010000e-07 V_low
+ 9.795000000e-07 V_low
+ 9.795010000e-07 V_low
+ 9.796000000e-07 V_low
+ 9.796010000e-07 V_low
+ 9.797000000e-07 V_low
+ 9.797010000e-07 V_low
+ 9.798000000e-07 V_low
+ 9.798010000e-07 V_low
+ 9.799000000e-07 V_low
+ 9.799010000e-07 V_hig
+ 9.800000000e-07 V_hig
+ 9.800010000e-07 V_hig
+ 9.801000000e-07 V_hig
+ 9.801010000e-07 V_hig
+ 9.802000000e-07 V_hig
+ 9.802010000e-07 V_hig
+ 9.803000000e-07 V_hig
+ 9.803010000e-07 V_hig
+ 9.804000000e-07 V_hig
+ 9.804010000e-07 V_hig
+ 9.805000000e-07 V_hig
+ 9.805010000e-07 V_hig
+ 9.806000000e-07 V_hig
+ 9.806010000e-07 V_hig
+ 9.807000000e-07 V_hig
+ 9.807010000e-07 V_hig
+ 9.808000000e-07 V_hig
+ 9.808010000e-07 V_hig
+ 9.809000000e-07 V_hig
+ 9.809010000e-07 V_hig
+ 9.810000000e-07 V_hig
+ 9.810010000e-07 V_hig
+ 9.811000000e-07 V_hig
+ 9.811010000e-07 V_hig
+ 9.812000000e-07 V_hig
+ 9.812010000e-07 V_hig
+ 9.813000000e-07 V_hig
+ 9.813010000e-07 V_hig
+ 9.814000000e-07 V_hig
+ 9.814010000e-07 V_hig
+ 9.815000000e-07 V_hig
+ 9.815010000e-07 V_hig
+ 9.816000000e-07 V_hig
+ 9.816010000e-07 V_hig
+ 9.817000000e-07 V_hig
+ 9.817010000e-07 V_hig
+ 9.818000000e-07 V_hig
+ 9.818010000e-07 V_hig
+ 9.819000000e-07 V_hig
+ 9.819010000e-07 V_hig
+ 9.820000000e-07 V_hig
+ 9.820010000e-07 V_hig
+ 9.821000000e-07 V_hig
+ 9.821010000e-07 V_hig
+ 9.822000000e-07 V_hig
+ 9.822010000e-07 V_hig
+ 9.823000000e-07 V_hig
+ 9.823010000e-07 V_hig
+ 9.824000000e-07 V_hig
+ 9.824010000e-07 V_hig
+ 9.825000000e-07 V_hig
+ 9.825010000e-07 V_hig
+ 9.826000000e-07 V_hig
+ 9.826010000e-07 V_hig
+ 9.827000000e-07 V_hig
+ 9.827010000e-07 V_hig
+ 9.828000000e-07 V_hig
+ 9.828010000e-07 V_hig
+ 9.829000000e-07 V_hig
+ 9.829010000e-07 V_low
+ 9.830000000e-07 V_low
+ 9.830010000e-07 V_low
+ 9.831000000e-07 V_low
+ 9.831010000e-07 V_low
+ 9.832000000e-07 V_low
+ 9.832010000e-07 V_low
+ 9.833000000e-07 V_low
+ 9.833010000e-07 V_low
+ 9.834000000e-07 V_low
+ 9.834010000e-07 V_low
+ 9.835000000e-07 V_low
+ 9.835010000e-07 V_low
+ 9.836000000e-07 V_low
+ 9.836010000e-07 V_low
+ 9.837000000e-07 V_low
+ 9.837010000e-07 V_low
+ 9.838000000e-07 V_low
+ 9.838010000e-07 V_low
+ 9.839000000e-07 V_low
+ 9.839010000e-07 V_hig
+ 9.840000000e-07 V_hig
+ 9.840010000e-07 V_hig
+ 9.841000000e-07 V_hig
+ 9.841010000e-07 V_hig
+ 9.842000000e-07 V_hig
+ 9.842010000e-07 V_hig
+ 9.843000000e-07 V_hig
+ 9.843010000e-07 V_hig
+ 9.844000000e-07 V_hig
+ 9.844010000e-07 V_hig
+ 9.845000000e-07 V_hig
+ 9.845010000e-07 V_hig
+ 9.846000000e-07 V_hig
+ 9.846010000e-07 V_hig
+ 9.847000000e-07 V_hig
+ 9.847010000e-07 V_hig
+ 9.848000000e-07 V_hig
+ 9.848010000e-07 V_hig
+ 9.849000000e-07 V_hig
+ 9.849010000e-07 V_hig
+ 9.850000000e-07 V_hig
+ 9.850010000e-07 V_hig
+ 9.851000000e-07 V_hig
+ 9.851010000e-07 V_hig
+ 9.852000000e-07 V_hig
+ 9.852010000e-07 V_hig
+ 9.853000000e-07 V_hig
+ 9.853010000e-07 V_hig
+ 9.854000000e-07 V_hig
+ 9.854010000e-07 V_hig
+ 9.855000000e-07 V_hig
+ 9.855010000e-07 V_hig
+ 9.856000000e-07 V_hig
+ 9.856010000e-07 V_hig
+ 9.857000000e-07 V_hig
+ 9.857010000e-07 V_hig
+ 9.858000000e-07 V_hig
+ 9.858010000e-07 V_hig
+ 9.859000000e-07 V_hig
+ 9.859010000e-07 V_hig
+ 9.860000000e-07 V_hig
+ 9.860010000e-07 V_hig
+ 9.861000000e-07 V_hig
+ 9.861010000e-07 V_hig
+ 9.862000000e-07 V_hig
+ 9.862010000e-07 V_hig
+ 9.863000000e-07 V_hig
+ 9.863010000e-07 V_hig
+ 9.864000000e-07 V_hig
+ 9.864010000e-07 V_hig
+ 9.865000000e-07 V_hig
+ 9.865010000e-07 V_hig
+ 9.866000000e-07 V_hig
+ 9.866010000e-07 V_hig
+ 9.867000000e-07 V_hig
+ 9.867010000e-07 V_hig
+ 9.868000000e-07 V_hig
+ 9.868010000e-07 V_hig
+ 9.869000000e-07 V_hig
+ 9.869010000e-07 V_low
+ 9.870000000e-07 V_low
+ 9.870010000e-07 V_low
+ 9.871000000e-07 V_low
+ 9.871010000e-07 V_low
+ 9.872000000e-07 V_low
+ 9.872010000e-07 V_low
+ 9.873000000e-07 V_low
+ 9.873010000e-07 V_low
+ 9.874000000e-07 V_low
+ 9.874010000e-07 V_low
+ 9.875000000e-07 V_low
+ 9.875010000e-07 V_low
+ 9.876000000e-07 V_low
+ 9.876010000e-07 V_low
+ 9.877000000e-07 V_low
+ 9.877010000e-07 V_low
+ 9.878000000e-07 V_low
+ 9.878010000e-07 V_low
+ 9.879000000e-07 V_low
+ 9.879010000e-07 V_hig
+ 9.880000000e-07 V_hig
+ 9.880010000e-07 V_hig
+ 9.881000000e-07 V_hig
+ 9.881010000e-07 V_hig
+ 9.882000000e-07 V_hig
+ 9.882010000e-07 V_hig
+ 9.883000000e-07 V_hig
+ 9.883010000e-07 V_hig
+ 9.884000000e-07 V_hig
+ 9.884010000e-07 V_hig
+ 9.885000000e-07 V_hig
+ 9.885010000e-07 V_hig
+ 9.886000000e-07 V_hig
+ 9.886010000e-07 V_hig
+ 9.887000000e-07 V_hig
+ 9.887010000e-07 V_hig
+ 9.888000000e-07 V_hig
+ 9.888010000e-07 V_hig
+ 9.889000000e-07 V_hig
+ 9.889010000e-07 V_hig
+ 9.890000000e-07 V_hig
+ 9.890010000e-07 V_hig
+ 9.891000000e-07 V_hig
+ 9.891010000e-07 V_hig
+ 9.892000000e-07 V_hig
+ 9.892010000e-07 V_hig
+ 9.893000000e-07 V_hig
+ 9.893010000e-07 V_hig
+ 9.894000000e-07 V_hig
+ 9.894010000e-07 V_hig
+ 9.895000000e-07 V_hig
+ 9.895010000e-07 V_hig
+ 9.896000000e-07 V_hig
+ 9.896010000e-07 V_hig
+ 9.897000000e-07 V_hig
+ 9.897010000e-07 V_hig
+ 9.898000000e-07 V_hig
+ 9.898010000e-07 V_hig
+ 9.899000000e-07 V_hig
+ 9.899010000e-07 V_hig
+ 9.900000000e-07 V_hig
+ 9.900010000e-07 V_hig
+ 9.901000000e-07 V_hig
+ 9.901010000e-07 V_hig
+ 9.902000000e-07 V_hig
+ 9.902010000e-07 V_hig
+ 9.903000000e-07 V_hig
+ 9.903010000e-07 V_hig
+ 9.904000000e-07 V_hig
+ 9.904010000e-07 V_hig
+ 9.905000000e-07 V_hig
+ 9.905010000e-07 V_hig
+ 9.906000000e-07 V_hig
+ 9.906010000e-07 V_hig
+ 9.907000000e-07 V_hig
+ 9.907010000e-07 V_hig
+ 9.908000000e-07 V_hig
+ 9.908010000e-07 V_hig
+ 9.909000000e-07 V_hig
+ 9.909010000e-07 V_low
+ 9.910000000e-07 V_low
+ 9.910010000e-07 V_low
+ 9.911000000e-07 V_low
+ 9.911010000e-07 V_low
+ 9.912000000e-07 V_low
+ 9.912010000e-07 V_low
+ 9.913000000e-07 V_low
+ 9.913010000e-07 V_low
+ 9.914000000e-07 V_low
+ 9.914010000e-07 V_low
+ 9.915000000e-07 V_low
+ 9.915010000e-07 V_low
+ 9.916000000e-07 V_low
+ 9.916010000e-07 V_low
+ 9.917000000e-07 V_low
+ 9.917010000e-07 V_low
+ 9.918000000e-07 V_low
+ 9.918010000e-07 V_low
+ 9.919000000e-07 V_low
+ 9.919010000e-07 V_low
+ 9.920000000e-07 V_low
+ 9.920010000e-07 V_low
+ 9.921000000e-07 V_low
+ 9.921010000e-07 V_low
+ 9.922000000e-07 V_low
+ 9.922010000e-07 V_low
+ 9.923000000e-07 V_low
+ 9.923010000e-07 V_low
+ 9.924000000e-07 V_low
+ 9.924010000e-07 V_low
+ 9.925000000e-07 V_low
+ 9.925010000e-07 V_low
+ 9.926000000e-07 V_low
+ 9.926010000e-07 V_low
+ 9.927000000e-07 V_low
+ 9.927010000e-07 V_low
+ 9.928000000e-07 V_low
+ 9.928010000e-07 V_low
+ 9.929000000e-07 V_low
+ 9.929010000e-07 V_hig
+ 9.930000000e-07 V_hig
+ 9.930010000e-07 V_hig
+ 9.931000000e-07 V_hig
+ 9.931010000e-07 V_hig
+ 9.932000000e-07 V_hig
+ 9.932010000e-07 V_hig
+ 9.933000000e-07 V_hig
+ 9.933010000e-07 V_hig
+ 9.934000000e-07 V_hig
+ 9.934010000e-07 V_hig
+ 9.935000000e-07 V_hig
+ 9.935010000e-07 V_hig
+ 9.936000000e-07 V_hig
+ 9.936010000e-07 V_hig
+ 9.937000000e-07 V_hig
+ 9.937010000e-07 V_hig
+ 9.938000000e-07 V_hig
+ 9.938010000e-07 V_hig
+ 9.939000000e-07 V_hig
+ 9.939010000e-07 V_hig
+ 9.940000000e-07 V_hig
+ 9.940010000e-07 V_hig
+ 9.941000000e-07 V_hig
+ 9.941010000e-07 V_hig
+ 9.942000000e-07 V_hig
+ 9.942010000e-07 V_hig
+ 9.943000000e-07 V_hig
+ 9.943010000e-07 V_hig
+ 9.944000000e-07 V_hig
+ 9.944010000e-07 V_hig
+ 9.945000000e-07 V_hig
+ 9.945010000e-07 V_hig
+ 9.946000000e-07 V_hig
+ 9.946010000e-07 V_hig
+ 9.947000000e-07 V_hig
+ 9.947010000e-07 V_hig
+ 9.948000000e-07 V_hig
+ 9.948010000e-07 V_hig
+ 9.949000000e-07 V_hig
+ 9.949010000e-07 V_low
+ 9.950000000e-07 V_low
+ 9.950010000e-07 V_low
+ 9.951000000e-07 V_low
+ 9.951010000e-07 V_low
+ 9.952000000e-07 V_low
+ 9.952010000e-07 V_low
+ 9.953000000e-07 V_low
+ 9.953010000e-07 V_low
+ 9.954000000e-07 V_low
+ 9.954010000e-07 V_low
+ 9.955000000e-07 V_low
+ 9.955010000e-07 V_low
+ 9.956000000e-07 V_low
+ 9.956010000e-07 V_low
+ 9.957000000e-07 V_low
+ 9.957010000e-07 V_low
+ 9.958000000e-07 V_low
+ 9.958010000e-07 V_low
+ 9.959000000e-07 V_low
+ 9.959010000e-07 V_hig
+ 9.960000000e-07 V_hig
+ 9.960010000e-07 V_hig
+ 9.961000000e-07 V_hig
+ 9.961010000e-07 V_hig
+ 9.962000000e-07 V_hig
+ 9.962010000e-07 V_hig
+ 9.963000000e-07 V_hig
+ 9.963010000e-07 V_hig
+ 9.964000000e-07 V_hig
+ 9.964010000e-07 V_hig
+ 9.965000000e-07 V_hig
+ 9.965010000e-07 V_hig
+ 9.966000000e-07 V_hig
+ 9.966010000e-07 V_hig
+ 9.967000000e-07 V_hig
+ 9.967010000e-07 V_hig
+ 9.968000000e-07 V_hig
+ 9.968010000e-07 V_hig
+ 9.969000000e-07 V_hig
+ 9.969010000e-07 V_low
+ 9.970000000e-07 V_low
+ 9.970010000e-07 V_low
+ 9.971000000e-07 V_low
+ 9.971010000e-07 V_low
+ 9.972000000e-07 V_low
+ 9.972010000e-07 V_low
+ 9.973000000e-07 V_low
+ 9.973010000e-07 V_low
+ 9.974000000e-07 V_low
+ 9.974010000e-07 V_low
+ 9.975000000e-07 V_low
+ 9.975010000e-07 V_low
+ 9.976000000e-07 V_low
+ 9.976010000e-07 V_low
+ 9.977000000e-07 V_low
+ 9.977010000e-07 V_low
+ 9.978000000e-07 V_low
+ 9.978010000e-07 V_low
+ 9.979000000e-07 V_low
+ 9.979010000e-07 V_hig
+ 9.980000000e-07 V_hig
+ 9.980010000e-07 V_hig
+ 9.981000000e-07 V_hig
+ 9.981010000e-07 V_hig
+ 9.982000000e-07 V_hig
+ 9.982010000e-07 V_hig
+ 9.983000000e-07 V_hig
+ 9.983010000e-07 V_hig
+ 9.984000000e-07 V_hig
+ 9.984010000e-07 V_hig
+ 9.985000000e-07 V_hig
+ 9.985010000e-07 V_hig
+ 9.986000000e-07 V_hig
+ 9.986010000e-07 V_hig
+ 9.987000000e-07 V_hig
+ 9.987010000e-07 V_hig
+ 9.988000000e-07 V_hig
+ 9.988010000e-07 V_hig
+ 9.989000000e-07 V_hig
+ 9.989010000e-07 V_hig
+ 9.990000000e-07 V_hig
+ 9.990010000e-07 V_hig
+ 9.991000000e-07 V_hig
+ 9.991010000e-07 V_hig
+ 9.992000000e-07 V_hig
+ 9.992010000e-07 V_hig
+ 9.993000000e-07 V_hig
+ 9.993010000e-07 V_hig
+ 9.994000000e-07 V_hig
+ 9.994010000e-07 V_hig
+ 9.995000000e-07 V_hig
+ 9.995010000e-07 V_hig
+ 9.996000000e-07 V_hig
+ 9.996010000e-07 V_hig
+ 9.997000000e-07 V_hig
+ 9.997010000e-07 V_hig
+ 9.998000000e-07 V_hig
+ 9.998010000e-07 V_hig
+ 9.999000000e-07 V_hig
+ 9.999010000e-07 V_hig
+ 1.000000000e-06 V_hig
+ 1.000001000e-06 V_hig
+ 1.000100000e-06 V_hig
+ 1.000101000e-06 V_hig
+ 1.000200000e-06 V_hig
+ 1.000201000e-06 V_hig
+ 1.000300000e-06 V_hig
+ 1.000301000e-06 V_hig
+ 1.000400000e-06 V_hig
+ 1.000401000e-06 V_hig
+ 1.000500000e-06 V_hig
+ 1.000501000e-06 V_hig
+ 1.000600000e-06 V_hig
+ 1.000601000e-06 V_hig
+ 1.000700000e-06 V_hig
+ 1.000701000e-06 V_hig
+ 1.000800000e-06 V_hig
+ 1.000801000e-06 V_hig
+ 1.000900000e-06 V_hig
+ 
.END
